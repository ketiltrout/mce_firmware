library ieee;
use ieee.std_logic_1164.all;

package command_pack is
   
end command_pack;