-- Copyright (c) 2003 SCUBA-2 Project
--                  All Rights Reserved

--  THIS IS UNPUBLISHED PROPRIETARY SOURCE CODE OF THE SCUBA-2 Project
--  The copyright notice above does not evidence any
--  actual or intended publication of such source code.

--  SOURCE CODE IS PROVIDED "AS IS". ALL EXPRESS OR IMPLIED CONDITIONS,
--  REPRESENTATIONS, AND WARRANTIES, INCLUDING ANY IMPLIED WARRANT OF
--  MERCHANTABILITY, SATISFACTORY QUALITY, FITNESS FOR A PARTICULAR
--  PURPOSE, OR NON-INFRINGEMENT, ARE DISCLAIMED, EXCEPT TO THE EXTENT
--  THAT SUCH DISCLAIMERS ARE HELD TO BE LEGALLY INVALID.

-- For the purposes of this code the SCUBA-2 Project consists of the
-- following organisations.

-- UKATC, Royal Observatory, Blackford Hill Edinburgh EH9 3HJ
-- UBC,   University of British Columbia, Physics & Astronomy Department,
--        Vancouver BC, V6T 1Z1

-- 
--
-- <revision control keyword substitutions e.g. $Id: tb_card_id_test_wrapper.vhd,v 1.2 2004/03/24 05:56:52 erniel Exp $>
--
-- Project:	      SCUBA-2
-- Author:	       Jonathan Jacob
-- Organisation:  UBC
--
-- Description:
-- 
--
-- Revision history:
-- Feb. 3 2004   - Initial version      - JJ
-- <date $Date: 2004/03/24 05:56:52 $>	-		<text>		- <initials $Author: erniel $>
-- $Log: tb_card_id_test_wrapper.vhd,v $
-- Revision 1.2  2004/03/24 05:56:52  erniel
-- added 8 more transmits
--
--
-----------------------------------------------------------------------------


library IEEE;
use IEEE.std_logic_1164.all;

library components;
use components.component_pack.all;

library sys_param;
use sys_param.wishbone_pack.all;


entity TB_CARD_ID_TEST_WRAPPER is
end TB_CARD_ID_TEST_WRAPPER;

architecture BEH of TB_CARD_ID_TEST_WRAPPER is

   component CARD_ID_TEST_WRAPPER
      port(RST_I       : in std_logic ;
           CLK_I       : in std_logic ;
           EN_I        : in std_logic ;
           DONE_O      : out std_logic ;
           TX_BUSY_I   : in std_logic ;
           TX_ACK_I    : in std_logic ;
           TX_DATA_O   : out std_logic_vector ( 7 downto 0 );
           TX_WE_O     : out std_logic ;
           TX_STB_O    : out std_logic ;
           DATA_BI     : inout std_logic );

   end component;


   constant PERIOD : time := 20 ns;

   signal W_RST_I       : std_logic ;
   signal W_CLK_I       : std_logic := '0';
   signal W_EN_I        : std_logic ;
   signal W_DONE_O      : std_logic ;
   signal W_TX_BUSY_I   : std_logic ;
   signal W_TX_ACK_I    : std_logic ;
   signal W_TX_DATA_O   : std_logic_vector ( 7 downto 0 );
   signal W_TX_WE_O     : std_logic ;
   signal W_TX_STB_O    : std_logic ;
   signal W_DATA_BI     : std_logic ;

   
   signal instr_command       : std_logic_vector(7 downto 0) := "00000000";

   constant SERIAL_CODE       : std_logic_vector(63 downto 0) :=  
                               "1000100011111111000000000000000011111111000000001111111100000000";
   -- alternate data for SERIAL_CODE:                           
   -- "0000111100001111000011110000111100001111000011110000111100001111";  -- 0x0F0F0F0F0F0F0F0F random data;
   -- "1000100011111111000000000000000011111111000000001111111100000000"   -- this is CRC calculated
   
   -- loop counters
   signal bit_count                    : integer := 1;
   signal i                            : integer := 8;
   
   -- reference data for self-checking
   signal reference_instr_command       : std_logic_vector(7 downto 0) := "00000000";
   signal reference_read_rom_cmd        : std_logic_vector(7 downto 0) := "00110011";
   

begin

------------------------------------------------------------------------
--
-- instantiate card_id_top
--
------------------------------------------------------------------------

   DUT : CARD_ID_TEST_WRAPPER
      port map(RST_I       => W_RST_I,
               CLK_I       => W_CLK_I,
               EN_I        => W_EN_I,
               DONE_O      => W_DONE_O,
               TX_BUSY_I   => W_TX_BUSY_I,
               TX_ACK_I    => W_TX_ACK_I,
               TX_DATA_O   => W_TX_DATA_O,
               TX_WE_O     => W_TX_WE_O,
               TX_STB_O    => W_TX_STB_O,
               DATA_BI     => W_DATA_BI);


------------------------------------------------------------------------
--
-- Create a test clock
--
------------------------------------------------------------------------

   W_CLK_I <= not W_CLK_I after PERIOD/2;
   
   

------------------------------------------------------------------------
--
-- Create stimulus
--
------------------------------------------------------------------------

   STIMULI : process
   
------------------------------------------------------------------------
--
-- Procdures for creating stimulus. MODEL THE ID CHIP, and the test interface
--
------------------------------------------------------------------------ 

      procedure do_nop is
      begin
      
         -- test software signals
         W_RST_I       <= '0';
         W_EN_I        <= '0';
         W_TX_BUSY_I   <= '0';
         W_TX_ACK_I    <= '0';
      
         -- ID chip signal
         W_DATA_BI   <= 'Z';
         
         wait for PERIOD;
         
         assert false report " Performing a NOP." severity NOTE;
      end do_nop ;
      
      
      procedure do_full_reset is
      begin
      
         -- test software signals
         W_RST_I       <= '1';
         W_EN_I        <= '0';
         W_TX_BUSY_I   <= '0';
         W_TX_ACK_I    <= '0';      
      
         -- ID chip signal
         W_DATA_BI   <= 'H';
         
         wait for PERIOD*3;

         -- test software signals
         W_RST_I       <= '0';
         W_EN_I        <= '0';
         W_TX_BUSY_I   <= '0';
         W_TX_ACK_I    <= '0';      
      
         -- ID chip signal
         W_DATA_BI   <= 'H';
         
         wait for PERIOD;
         
         assert false report " Performing a RESET." severity NOTE;
      end do_full_reset ;      


      procedure do_start is
      begin
      
         -- test software signals
         W_RST_I       <= '0';
         W_EN_I        <= '1';
         W_TX_BUSY_I   <= '0';
         W_TX_ACK_I    <= '0';   

         -- ID chip pulling bus high
         W_DATA_BI             <= 'H';
         
         wait for PERIOD;
         
         assert false report " STARTING the TEST." severity NOTE;
      end do_start ;     



      procedure do_id_chip_init_pulse is
         begin
      
         W_DATA_BI             <= 'H';    
         wait for 400 us;
      
         wait until W_DATA_BI  <= 'H';
         
         -- this is the ID chip pulling the bus low
         wait for 15 us;
         W_DATA_BI             <= '0';
         wait for 60 us;
         -- release the bus
         W_DATA_BI             <= 'H';
      
         wait for PERIOD;

         assert false report "Presence Pulse is done";
      end do_id_chip_init_pulse;


      procedure do_id_chip_read_rom_cmd is
      begin
      
      while i > 0 loop

         W_DATA_BI   <= 'H';
        
         assert false report " Master is writing 0x33 to the DS18S20 " severity NOTE;

         wait until W_DATA_BI   <= '0';

         wait for 40 us;   
         
         -- sample the data and shift it into instr_command register
         instr_command <= W_DATA_BI & instr_command(7 downto 1);
         
         -- this is the reference data for the self-checking
         reference_instr_command <= reference_read_rom_cmd(8-i) & reference_instr_command(7 downto 1);
         
         i <= i-1;       
         wait for 20 us;
         
         -- self-checking: bit pattern during shift in should be
         -- 10000000 0x80 shift 1
         -- 11000000 0xC0 shift 2
         -- 01100000 0x60 shift 3
         -- 00110000 0x30 shift 4
         -- 10110000 0xB0 shift 5
         -- 11001100 0xCC shift 6
         -- 01100110 0x66 shift 7
         -- 00110011 0x33 shift 8
        
         --assert instr_command = reference_instr_command report " SELF-CHECKING FAILED DURING 'READ ROM' COMMAND " severity FAILURE;
      
        end loop; 
     end do_id_chip_read_rom_cmd; 
   

     procedure do_master_sample is
     begin
      
         while bit_count < 64 loop

         wait until W_DATA_BI = '0';

         wait for 4 us;   
         
         -- Output the family code, serial code and CRC one bit at a time
         -- This is the data coming from the ID chip
         if SERIAL_CODE(bit_count-1) = '1' then
            W_DATA_BI <= 'H';
         else
            W_DATA_BI <= 'L';
         end if;   
         assert false report " Master is sampling bit from the DS18S20 " severity NOTE;
        
         wait for 56 us;
         bit_count <= bit_count + 1;     
         W_DATA_BI                 <= 'H';        
                  
         end loop;
         
      end do_master_sample; 


      procedure do_wait is
      begin
      
         wait for PERIOD;
         
         -- test software signals
         W_RST_I       <= '0';
         W_EN_I        <= '1';
         W_TX_BUSY_I   <= '0';
         W_TX_ACK_I    <= '0';      
      
         -- ID chip signal
         W_DATA_BI   <= 'H';      

         wait for 10 us;        
         
         assert false report " Waiting for 10 us." severity NOTE;
      end do_wait ;     
      
 
 
      procedure do_tx_byte_to_RS232 is
      begin


         -- this means the test wrapper is ready to send data to the RS232
         if w_tx_stb_o = '0' then
            wait until w_tx_stb_o = '1';
         end if;
         
         if w_tx_we_o = '0' then
            wait until w_tx_we_o = '1';
         end if;
         
         -- test software signals
         W_RST_I       <= '0';
         W_EN_I        <= '1';
         W_TX_BUSY_I   <= '0';
         W_TX_ACK_I    <= '1';  -- grab the data
         
         wait for PERIOD;
         
         W_RST_I       <= '0';
         W_EN_I        <= '1';
         W_TX_BUSY_I   <= '1';  -- indicates it's busy now writing the "grabbed" data to the RS232
         W_TX_ACK_I    <= '0';
         
         
         wait for PERIOD*3;
         
         W_RST_I       <= '0';
         W_EN_I        <= '1';
         W_TX_BUSY_I   <= '0';
         W_TX_ACK_I    <= '0';   
         
         wait for PERIOD;      
         
         assert false report " Writing out the data to RS232." severity NOTE;
      end do_tx_byte_to_RS232;    


      procedure do_tx_byte_to_RS232_last is
      begin


         -- this means the test wrapper is ready to send data to the RS232
         if w_tx_stb_o = '0' then
            wait until w_tx_stb_o = '1';
         end if;
         
         if w_tx_we_o = '0' then
            wait until w_tx_we_o = '1';
         end if;
         
         -- test software signals
         W_RST_I       <= '0';
         W_EN_I        <= '1';
         W_TX_BUSY_I   <= '0';
         W_TX_ACK_I    <= '1';  -- grab the data
         
         wait until w_done_o = '0';
         
         W_RST_I       <= '0';
         W_EN_I        <= '0';
         W_TX_BUSY_I   <= '1';  -- indicates it's busy now writing the "grabbed" data to the RS232
         W_TX_ACK_I    <= '0';
         
         
         wait for PERIOD*3;
         
         W_RST_I       <= '0';
         W_EN_I        <= '0';
         W_TX_BUSY_I   <= '0';
         W_TX_ACK_I    <= '0';   
         
         wait for PERIOD;  
         
         assert false report " Writing out the data to RS232." severity NOTE;
      end do_tx_byte_to_RS232_last;  




      procedure do_finish is
      begin
      
         wait until W_DONE_O = '1';

         wait for PERIOD;
         
         -- test software signals
         W_RST_I       <= '0';
         W_EN_I        <= '0';
         W_TX_BUSY_I   <= '0';
         W_TX_ACK_I    <= '0';      
      
         -- ID chip signal
         W_DATA_BI   <= 'H';      

         wait for 10 us;     
 
         assert false report " Finishing up..." severity NOTE;
      end do_finish ;     

------------------------------------------------------------------------
--
-- Start the test
--
------------------------------------------------------------------------
          
   begin
      do_nop;
      
      do_full_reset;  
      
      do_start;
      

      do_id_chip_init_pulse;
      
      do_id_chip_read_rom_cmd;
      
      do_master_sample;
             
      do_wait;

      do_tx_byte_to_RS232;
      do_tx_byte_to_RS232;
      do_tx_byte_to_RS232;
      do_tx_byte_to_RS232;
      
      do_tx_byte_to_RS232;
      do_tx_byte_to_RS232;
      do_tx_byte_to_RS232;
      do_tx_byte_to_RS232;
      
      do_tx_byte_to_RS232;
      do_tx_byte_to_RS232;
      do_tx_byte_to_RS232;
      do_tx_byte_to_RS232;
      
      do_tx_byte_to_RS232;
      do_tx_byte_to_RS232;
      do_tx_byte_to_RS232;
      do_tx_byte_to_RS232;
      
--      do_tx_byte_to_RS232_last;

      do_finish;
      
      assert false report " FINISHED: Simulation done." severity FAILURE;
      
   end process STIMULI;

end beh;
