-- Copyright (c) 2003 SCUBA-2 Project
-- All Rights Reserved
--
-- THIS IS UNPUBLISHED PROPRIETARY SOURCE CODE OF THE SCUBA-2 Project
-- The copyright notice above does not evidence any
-- actual or intended publication of such source code.
--
-- SOURCE CODE IS PROVIDED "AS IS". ALL EXPRESS OR IMPLIED CONDITIONS,
-- REPRESENTATIONS, AND WARRANTIES, INCLUDING ANY IMPLIED WARRANT OF
-- MERCHANTABILITY, SATISFACTORY QUALITY, FITNESS FOR A PARTICULAR
-- PURPOSE, OR NON-INFRINGEMENT, ARE DISCLAIMED, EXCEPT TO THE EXTENT
-- THAT SUCH DISCLAIMERS ARE HELD TO BE LEGALLY INVALID.
--
-- For the purposes of this code the SCUBA-2 Project consists of the
-- following organisations.
--
-- UKATC, Royal Observatory, Blackford Hill Edinburgh EH9 3HJ
-- UBC, University of British Columbia, Physics & Astronomy Department,
-- Vancouver BC, V6T 1Z1
--
-- tb_tx_reply
--
--
-- Project: 			Scuba 2
-- Author:  			David Atkinson
-- Organisation: 			UKATC
--
-- Description:
-- test bed for tx_reply
--
-- Revision history:
-- <date $Date: 2004/10/08 14:10:32 $> - <text> - <initials $Author: dca $>
--
-- $Log: tb_tx_reply.vhd,v $
-- Revision 1.1  2004/10/08 14:10:32  dca
-- Initial version
--
--
-- 
-----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity tb_tx_reply is
end tb_tx_reply;



library ieee;
use ieee.std_logic_1164.all;

library work;
use work.issue_reply_pack.all;

library sys_param;
use sys_param.command_pack.all;
use sys_param.wishbone_pack.all;


architecture bench of tb_tx_reply is


-- component declaration


------------------
component tx_reply
------------------
port(

-- global inputs 
   rst_i                   : in  std_logic;                                            -- global reset
   clk_i                   : in  std_logic;                                            -- global clock

-- signals to/from cmd_translator    
   cmd_rcvd_er_i           : in  std_logic;                                            -- command received on fibre with checksum error
   cmd_rcvd_ok_i           : in  std_logic;                                            -- command received on fibre - no checksum error
   cmd_code_i              : in  std_logic_vector (FIBRE_CMD_CODE_WIDTH-1  downto 0);    -- fibre command code
   card_id_i               : in  std_logic_vector (FIBRE_CARD_ADDRESS_WIDTH-1 downto 0);    -- fibre command card id
   param_id_i              : in  std_logic_vector (FIBRE_PARAMETER_ID_WIDTH-1    downto 0);    -- fibre command parameter id
         
-- signals to/from reply queue 
   m_op_done_i             : in  std_logic;                                            -- macro op done
   m_op_ok_nEr_i           : in  std_logic;                                            -- macro op success ('1') or error ('0') 
   m_op_cmd_code_i         : in  std_logic_vector (BB_COMMAND_TYPE_WIDTH-1      downto 0);    -- command code vector - indicates if data or reply (and which command)
   fibre_word_i            : in  std_logic_vector (PACKET_WORD_WIDTH-1      downto 0);    -- packet word read from reply queue
   num_fibre_words_i       : in  std_logic_vector (PACKET_WORD_WIDTH-1      downto 0);    -- indicate number of packet words to be read from reply queue
   fibre_word_req_o        : out std_logic;                                            -- asserted to requeset next fibre word
   m_op_ack_o              : out std_logic;                                            -- asserted to indicate to reply queue the the packet has been processed

-- interface to HOTLINK transmitter
   ft_clkw_i               : in     std_logic;                                         -- HOTLINK clock - generated by FPGA
   nTrp_i                  : in     std_logic;                                         -- HOTLINK read pulse (to read tx FIFO)
   tx_data_o               : out    std_logic_vector(TX_FIFO_DATA_WIDTH-1 downto 0);   -- HOTLINK data byte to transmit
   tsc_nTd_o               : out    std_logic;                                         -- HOTLINK transmit special char / data select
   nFena_o                 : out    std_logic                                          -- HOTLINK transmit enable 
     );      
end component;


--------------------------
component tx_hotlink_sim
--------------------------
port( 
   ft_clkw_i              : in     std_logic;                                           -- HOTLINK clock - generated by FPGA
   nFena_i                : in     std_logic;                                           -- HOTLINK transmit enable 
   tsc_nTd_i              : in     std_logic;                                           -- HOTLINK transmit special char / data select  
   tx_data_i              : in     std_logic_vector (7 downto 0);                       -- HOTLINK data byte to transmit
   nTrp_o                 : out    std_logic                                            -- HOTLINK read pulse (to read tx FIFO)
   );
end component;


-- signal declarations


-- signals to/from cmd_translator    
signal    cmd_rcvd_er        : std_logic := '0';                                                      -- command received on fibre with checksum error
signal    cmd_rcvd_ok        : std_logic := '0';                                                      -- command received on fibre - no checksum error
signal    cmd_code           : std_logic_vector (FIBRE_CMD_CODE_WIDTH-1  downto 0) := (others => '0');  -- fibre command code
signal    card_id            : std_logic_vector (FIBRE_CARD_ADDRESS_WIDTH-1 downto 0) := (others => '0');  -- fibre command card id
signal    param_id           : std_logic_vector (FIBRE_PARAMETER_ID_WIDTH-1    downto 0) := (others => '0');  -- fibre command parameter id
         
-- signals to/from reply queue 
signal    m_op_done          : std_logic;                                             -- macro op done
signal    m_op_ok_nEr        : std_logic;                                             -- macro op success ('1') or error ('0') 
signal    m_op_cmd_code      : std_logic_vector (BB_COMMAND_TYPE_WIDTH-1      downto 0);     -- command code vector - indicates if data or reply (and which command)
signal    fibre_word         : std_logic_vector (PACKET_WORD_WIDTH-1      downto 0);     -- packet word read from reply queue
signal    num_fibre_words    : std_logic_vector (PACKET_WORD_WIDTH-1      downto 0);     -- indicate number of packet words to be read from reply queue
signal    fibre_word_req     : std_logic;                                             -- asserted to requeset next fibre word
signal    m_op_ack           : std_logic;                                             -- asserted to indicate to reply queue the the packet has been processed

-- interface to HOTLINK transmitter
signal   ft_clkw             : std_logic := '0';                                  -- HOTLINK clock - generated by FPGA
signal   nTrp                : std_logic;                                         -- HOTLINK read pulse (to read tx FIFO)
signal   tx_data             : std_logic_vector(TX_FIFO_DATA_WIDTH-1 downto 0);   -- HOTLINK data byte to transmit
signal   tsc_nTd             : std_logic;                                         -- HOTLINK transmit special char / data select
signal   nFena               : std_logic;                                         -- HOTLINK transmit enable 

signal   tb_clk              : std_logic := '0';
signal   dut_rst             : std_logic;
           
constant clk_prd      : TIME := 20 ns;    -- 50Mhz clock 
constant ft_clkw_prd  : TIME := 40 ns;    -- 25Mhz clock
 
begin

   -- Instantiate design under test
   DUT : tx_reply
   port map(

   -- global inputs 
      rst_i             =>  dut_rst, 
      clk_i             =>  tb_clk,

   -- signals to/from cmd_translator    
      cmd_rcvd_er_i     =>  cmd_rcvd_er,                                   
      cmd_rcvd_ok_i     =>  cmd_rcvd_ok,
      cmd_code_i        =>  cmd_code,
      card_id_i         =>  card_id,
      param_id_i        =>  param_id,
         
   -- signals to/from reply queue 
      m_op_done_i       =>  m_op_done,
      m_op_ok_nEr_i     =>  m_op_ok_nEr,                                         
      m_op_cmd_code_i   =>  m_op_cmd_code,
      fibre_word_i      =>  fibre_word,
      num_fibre_words_i =>  num_fibre_words,
      fibre_word_req_o  =>  fibre_word_req,
      m_op_ack_o        =>  m_op_ack,

   -- interface to HOTLINK transmitter
      ft_clkw_i         =>  ft_clkw,
      nTrp_i            =>  nTrp,
      tx_data_o         =>  tx_data,
      tsc_nTd_o         =>  tsc_nTd,
      nFena_o           =>  nFena
     );      
   
   -- instantiate holink transmitter simulator
   
   SIM : tx_hotlink_sim
   port map(
   
      ft_clkw_i         =>  ft_clkw,
      nFena_i           =>  nFena,
      tsc_nTd_i         =>  tsc_nTd,  
      tx_data_i         =>  tx_data,
      nTrp_o            =>  nTrp
   );
           
         
------------------------------------------------
-- Create test bench clock
-------------------------------------------------
  
   tb_clk <= not tb_clk after clk_prd/2;

        
------------------------------------------------
-- Create hotlink sim clock 
-------------------------------------------------
  
   ft_clkw <= not ft_clkw after ft_clkw_prd/2;
   
------------------------------------------------
-- Create test bench stimuli
-------------------------------------------------
   
   stimuli : process
  
------------------------------------------------
-- Stimulus procedures
-------------------------------------------------
      
   procedure do_reset is
   begin
      dut_rst <= '1';
      assert false report " Resetting the DUT." severity NOTE;
      wait for clk_prd*5 ;
      dut_rst <= '0';
      wait for clk_prd*5 ;
   
      
   end do_reset;
--------------------------------------------------         
   
   begin 
      dut_rst <= '0';
      wait for clk_prd*5;
      
      do_reset;
      
      -- generate a checksum error reply
      cmd_code      <= ASCII_R & ASCII_B;
      card_id       <= X"0012";
      param_id      <= X"010C";
      cmd_rcvd_er   <= '1'; 
      wait for clk_prd*5;
      cmd_rcvd_er  <= '0';
      wait for clk_prd*5;
      
      
      for i in 1 to 30 loop
         wait until nTrp = '0';
         assert false report "Byte Requested" severity NOTE;
      end loop;
      
      wait for clk_prd*30;
 
      assert false report "Simulation done." severity FAILURE;
      wait ;

   end process stimuli;         
           
end bench;