-- Copyright (c) 2003 SCUBA-2 Project
--                  All Rights Reserved

--  THIS IS UNPUBLISHED PROPRIETARY SOURCE CODE OF THE SCUBA-2 Project
--  The copyright notice above does not evidence any
--  actual or intended publication of such source code.

--  SOURCE CODE IS PROVIDED "AS IS". ALL EXPRESS OR IMPLIED CONDITIONS,
--  REPRESENTATIONS, AND WARRANTIES, INCLUDING ANY IMPLIED WARRANT OF
--  MERCHANTABILITY, SATISFACTORY QUALITY, FITNESS FOR A PARTICULAR
--  PURPOSE, OR NON-INFRINGEMENT, ARE DISCLAIMED, EXCEPT TO THE EXTENT
--  THAT SUCH DISCLAIMERS ARE HELD TO BE LEGALLY INVALID.

-- For the purposes of this code the SCUBA-2 Project consists of the
-- following organisations.

-- UKATC, Royal Observatory, Blackford Hill Edinburgh EH9 3HJ
-- UBC,   University of British Columbia, Physics & Astronomy Department,
--        Vancouver BC, V6T 1Z1

-- frame_timing_pack.vhd
--
-- <revision control keyword substitutions e.g. $Id: frame_timing_pack.vhd,v 1.5 2004/05/14 21:10:06 mandana Exp $>
--
-- Project:     SCUBA-2
-- Author:      Bryce Burger
-- Organisation:  UBC
--
-- Description:
-- This records all of the constants needed for frame synchronization
-- on the AC, BC, RC.
--
-- Revision history:
-- <date $Date: 2004/05/14 21:10:06 $> - <text> - <initials $Author: mandana $>
-- $Log: frame_timing_pack.vhd,v $
-- Revision 1.5  2004/05/14 21:10:06  mandana
-- changed frame_timing values to integer(Bias_count)
--
-- Revision 1.4  2004/05/13 00:09:10  bburger
-- added a few timing parameters for the clock card
--
-- Revision 1.3  2004/04/16 21:58:43  bburger
-- changed port names
--
-- Revision 1.2  2004/04/16 00:41:16  bburger
-- renamed some signals
--
-- Revision 1.1  2004/04/14 21:56:40  jjacob
-- new directory structure
--
-- Revision 1.6  2004/04/14 20:14:14  bburger
-- no message
--
-- Revision 1.5  2004/04/02 01:12:04  bburger
-- added a log field to header
--
--
------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

-- This package contains the timing information for the cards in the
-- MCE that need to be synchronized to an overall frame structure.
-- The frame structure is resolved to 50Mhz clock cycles.
-- If the resolution freqency changes, then all the constants below
-- will need to be adjusted.
-- Multiplexing by the MCE will occur at 781.250kHz, meaning that
-- address-dwell times will be 1.280us or the duration of 64 50MHz
-- cycles.
library sys_param;
use sys_param.data_types_pack.all;

package frame_timing_pack is

   constant MUX_LINE_PERIOD   : integer := 64; -- 64 50MHz cycles
   constant END_OF_FRAME      : integer := 41*MUX_LINE_PERIOD; --(41*MUX_LINE_PERIOD);

   ------------------------------------------------------------------------------------
   -- Clock Card frame structure

   -- START_OF_BLACKOUT:
   -- This value is used by the cmd_queue to determe whether it can issue a command.
   -- START_OF_BLACKOUT indicates the point in a frame at which there is not enough
   -- time remaining to send out a command and have the wishbone master parse it before
   -- data becomes invalid.
   -- During normal operation, there should be enough time in a frame to issue all
   -- required commands for normal operaiton.  However, START_OF_BLACKOUT may come
   -- into consideration if a corrupted reply was received by the reply_queue and
   -- the cmd_queue needs to reissued the corresponding u-op
   constant START_OF_BLACKOUT : integer := END_OF_FRAME - 5*MUX_LINE_PERIOD;

   -- RETIRE_TIMEOUT indicates at what point in a frame all the commands that were
   -- in that frame must be retired.
   -- If some commands remain to be retired at the end of a frame, some type of error
   -- recovery must be initiated
   constant RETIRE_TIMEOUT    : integer := END_OF_FRAME;

   ------------------------------------------------------------------------------------
   -- Bias Card frame structure
   constant UPDATE_BIAS : integer := 3;
   ------------------------------------------------------------------------------------
   -- Address Card frame structure
   constant SEL_ROW : w_array41:= (
    0*MUX_LINE_PERIOD,1*MUX_LINE_PERIOD, 2*MUX_LINE_PERIOD, 3*MUX_LINE_PERIOD, 4*MUX_LINE_PERIOD, 
    5*MUX_LINE_PERIOD, 6*MUX_LINE_PERIOD, 7*MUX_LINE_PERIOD, 8*MUX_LINE_PERIOD, 9*MUX_LINE_PERIOD,
    10*MUX_LINE_PERIOD,11*MUX_LINE_PERIOD,12*MUX_LINE_PERIOD,13*MUX_LINE_PERIOD,14*MUX_LINE_PERIOD,
    15*MUX_LINE_PERIOD,16*MUX_LINE_PERIOD,17*MUX_LINE_PERIOD,18*MUX_LINE_PERIOD,19*MUX_LINE_PERIOD,
    20*MUX_LINE_PERIOD,21*MUX_LINE_PERIOD,22*MUX_LINE_PERIOD,23*MUX_LINE_PERIOD,24*MUX_LINE_PERIOD,
    25*MUX_LINE_PERIOD,26*MUX_LINE_PERIOD,27*MUX_LINE_PERIOD,28*MUX_LINE_PERIOD,29*MUX_LINE_PERIOD,
    30*MUX_LINE_PERIOD,31*MUX_LINE_PERIOD,32*MUX_LINE_PERIOD,33*MUX_LINE_PERIOD,34*MUX_LINE_PERIOD,
    35*MUX_LINE_PERIOD,36*MUX_LINE_PERIOD,37*MUX_LINE_PERIOD,38*MUX_LINE_PERIOD,39*MUX_LINE_PERIOD, 
    40*MUX_LINE_PERIOD);

   ------------------------------------------------------------------------------------
   -- Frame Timing Interface

   component frame_timing is
   port(
         clk_i       : in std_logic;
         sync_i      : in std_logic;
         frame_rst_i : in std_logic;
         clk_count_o : out integer;
         clk_error_o : out std_logic_vector(31 downto 0)
      );
   end component;


end frame_timing_pack;