-- 2003 SCUBA-2 Project
--                  All Rights Reserved

--  THIS IS UNPUBLISHED PROPRIETARY SOURCE CODE OF THE SCUBA-2 Project
--  The copyright notice above does not evidence any
--  actual or intended publication of such source code.

--  SOURCE CODE IS PROVIDED "AS IS". ALL EXPRESS OR IMPLIED CONDITIONS,
--  REPRESENTATIONS, AND WARRANTIES, INCLUDING ANY IMPLIED WARRANT OF
--  MERCHANTABILITY, SATISFACTORY QUALITY, FITNESS FOR A PARTICULAR
--  PURPOSE, OR NON-INFRINGEMENT, ARE DISCLAIMED, EXCEPT TO THE EXTENT
--  THAT SUCH DISCLAIMERS ARE HELD TO BE LEGALLY INVALID.

-- For the purposes of this code the SCUBA-2 Project consists of the
-- following organisations.

-- UKATC, Royal Observatory, Blackford Hill Edinburgh EH9 3HJ
-- UBC,   University of British Columbia, Physics & Astronomy Department,
--        Vancouver BC, V6T 1Z1

-- $Id: bc_dac_ctrl.vhd,v 1.15 2016/05/19 22:12:19 mandana Exp $
--
-- Project:       SCUBA2
-- Author:        Bryce Burger
-- Organisation:  UBC
--
-- Description:
-- This block (and lower level blocks) processes wishbone commands and 
-- updates 32 flux_fb SPI DACs and 12 low-noise bias SPI DACs.
-- Wishbone commands processed by this block are:
-- FLUX_FB_ADDR 
-- BIAS_ADDR 
-- ENBL_MUX_ADDR
-- ENBL_FLUX_FB_MOD_ADDR
-- ENBL_BIAS_MOD_ADDR
-- MOD_VAL_ADDR
-- FB_COLxx
--
-- Revision history:
-- $Log: bc_dac_ctrl.vhd,v $
-- Revision 1.15  2016/05/19 22:12:19  mandana
-- 6.0.1 added flux_fb_dly parameter and removed num_idle_rows implementation
--
-- Revision 1.14  2014/12/18 23:21:41  mandana
-- 5.3.5 added num_idle_rows
--
-- Revision 1.13  2012-03-26 21:54:12  mandana
-- added comment about new commands!
--
-- Revision 1.12  2011-11-29 00:55:44  mandana
-- ln_bias_changed changed to std_logic_vector, one bit per DAC
--
-- Revision 1.11  2011-10-26 18:26:32  mandana
-- *** empty log message ***
--
-- Revision 1.10  2010/06/02 17:41:22  mandana
-- flux_fb_changed flag is now defined as 1 bit per column
-- 1row_prev is added to the interface
--
-- Revision 1.9  2010/05/14 00:03:24  mandana
-- added interface ports to read enbl_mux and mux_flux_fb_data
-- added ports for row_switch_i to the interface
--
-- Revision 1.8  2010/01/20 23:04:47  mandana
-- added interface for low-noise bias lines introduced in bias-card Rev. E
-- spi_clk_i or DAC clocks are now generated by PLL
--
-- Revision 1.7  2006/08/03 19:06:31  mandana
-- reorganized pack files, bc_dac_ctrl_core_pack, bc_dac_ctrl_wbs_pack, frame_timing_pack are all obsolete
--
-- Revision 1.6  2005/01/17 23:01:04  mandana
-- removed mem_clk_i
-- read from RAM is performed in 2 clk_i cycles, added an extra state for read
--
-- Revision 1.5  2005/01/04 19:19:47  bburger
-- Mandana: changed mictor assignment to 0 to 31 and swapped odd and even pods
--
-- Revision 1.4  2004/12/21 22:06:51  bburger
-- Bryce:  update
--
-- Revision 1.3  2004/11/25 03:05:08  bburger
-- Bryce:  Modified the Bias Card DAC control slaves.
--
-- Revision 1.2  2004/11/15 20:03:41  bburger
-- Bryce :  Moved frame_timing to the 'work' library, and physically moved the files to "all_cards" directory
--
-- Revision 1.1  2004/11/11 01:47:10  bburger
-- Bryce:  new
--
--   
--
-- 
-----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

library sys_param;
use sys_param.wishbone_pack.all;

library work;
use work.bias_card_pack.all;
use work.bc_dac_ctrl_pack.all;

entity bc_dac_ctrl is
   port
   (
      -- DAC hardware interface:
      -- 32 independant flux-fb DAC channels, thus 32 serial data/cs/clk lines and
      -- 12 ln_bias DAC channels, data and clk lines are shared
      flux_fb_data_o    : out std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);   
      flux_fb_ncs_o     : out std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);
      flux_fb_clk_o     : out std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);      
      
      ln_bias_data_o    : out std_logic;
      ln_bias_ncs_o     : out std_logic_vector(NUM_LN_BIAS_DACS-1 downto 0);
      ln_bias_clk_o     : out std_logic;
      
      dac_nclr_o        : out std_logic;
      
      -- wishbone interface:
      dat_i             : in std_logic_vector(WB_DATA_WIDTH-1 downto 0);
      addr_i            : in std_logic_vector(WB_ADDR_WIDTH-1 downto 0);
      tga_i             : in std_logic_vector(WB_TAG_ADDR_WIDTH-1 downto 0);
      we_i              : in std_logic;
      stb_i             : in std_logic;
      cyc_i             : in std_logic;
      dat_o             : out std_logic_vector(WB_DATA_WIDTH-1 downto 0);
      ack_o             : out std_logic;
      
      -- frame_timing signals
      row_switch_i      : in std_logic;
      update_bias_i     : in std_logic;
      flux_fb_dly_i     : in std_logic;
      restart_frame_aligned_i : in std_logic;      
      restart_frame_1row_prev_i : in std_logic;
      
      -- Global Signals      
      clk_i             : in std_logic;
      spi_clk_i         : in std_logic;
      rst_i             : in std_logic;
      debug             : inout std_logic_vector(31 downto 0)
   );     
end bc_dac_ctrl;

architecture rtl of bc_dac_ctrl is

   -- wbs_bc_dac_ctrl interface:
   signal flux_fb_addr    : std_logic_vector(FLUX_FB_DAC_ADDR_WIDTH-1 downto 0);
   signal flux_fb_data    : flux_fb_dac_array;--std_logic_vector(FLUX_FB_DAC_DATA_WIDTH-1 downto 0);
   signal flux_fb_changed : std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);
   signal ln_bias_addr    : std_logic_vector(LN_BIAS_DAC_ADDR_WIDTH-1 downto 0);
   signal ln_bias_data    : std_logic_vector(LN_BIAS_DAC_DATA_WIDTH-1 downto 0);
   signal ln_bias_changed : std_logic_vector(NUM_LN_BIAS_DACS-1 downto 0);   
   signal row_addr        : std_logic_vector(ROW_ADDR_WIDTH-1 downto 0);
   signal mux_flux_fb_data: flux_fb_dac_array;
   signal enbl_mux_data   : std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);
   
begin

   bcdc_core: bc_dac_ctrl_core
   port map(
      -- DAC hardware interface:
      flux_fb_data_o    => flux_fb_data_o,
      flux_fb_ncs_o     => flux_fb_ncs_o, 
      flux_fb_clk_o     => flux_fb_clk_o, 
      
      ln_bias_data_o    => ln_bias_data_o,
      ln_bias_ncs_o     => ln_bias_ncs_o, 
      ln_bias_clk_o     => ln_bias_clk_o, 
      
      dac_nclr_o        => dac_nclr_o,

      -- wbs_bc_dac_ctrl interface:
      row_addr_o        => row_addr,
      flux_fb_addr_o    => flux_fb_addr,
      flux_fb_data_i    => flux_fb_data,   
      flux_fb_changed_i => flux_fb_changed,
      ln_bias_addr_o    => ln_bias_addr,
      ln_bias_data_i    => ln_bias_data,      
      ln_bias_changed_i => ln_bias_changed,   

      mux_flux_fb_data_i=> mux_flux_fb_data,
      enbl_mux_data_i   => enbl_mux_data,
      
      -- frame_timing signals
      row_switch_i      => row_switch_i,
      update_bias_i     => update_bias_i,
      flux_fb_dly_i     => flux_fb_dly_i,
      restart_frame_aligned_i => restart_frame_aligned_i,
      restart_frame_1row_prev_i => restart_frame_1row_prev_i,

      -- Global Signals      
      clk_i             => clk_i,
      spi_clk_i         => spi_clk_i,
      rst_i             => rst_i,
      debug             => debug
   );     
       
   -- handles wishbone transactions  
   bcdc_wbs: bc_dac_ctrl_wbs
   port map(
      -- bc_dac_ctrl interface: 32 flux_fb DACs and up to 12 low-noise bias DACs
      flux_fb_addr_i    => flux_fb_addr,
      flux_fb_data_o    => flux_fb_data,   
      flux_fb_changed_o => flux_fb_changed,
      ln_bias_addr_i    => ln_bias_addr,
      ln_bias_data_o    => ln_bias_data,      
      ln_bias_changed_o => ln_bias_changed,   
     
      mux_flux_fb_data_o => mux_flux_fb_data,
      enbl_mux_data_o   => enbl_mux_data,
      row_addr_i        => row_addr,
      row_switch_i      => row_switch_i,
      
      -- wishbone interface:
      dat_i             => dat_i, 
      addr_i            => addr_i,
      tga_i             => tga_i, 
      we_i              => we_i,  
      stb_i             => stb_i, 
      cyc_i             => cyc_i, 
      dat_o             => dat_o, 
      ack_o             => ack_o, 

      -- global interface
      clk_i             => clk_i,
      rst_i             => rst_i,
      debug             => debug
   );
      
end rtl;