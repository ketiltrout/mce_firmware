-- megafunction wizard: %RAM: 3-PORT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: alt3pram 

-- ============================================================
-- File Name: cmd_queue_ram40.vhd
-- Megafunction Name(s):
-- 			alt3pram
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
-- ************************************************************


--Copyright (C) 1991-2003 Altera Corporation
--Any  megafunction  design,  and related netlist (encrypted  or  decrypted),
--support information,  device programming or simulation file,  and any other
--associated  documentation or information  provided by  Altera  or a partner
--under  Altera's   Megafunction   Partnership   Program  may  be  used  only
--to program  PLD  devices (but not masked  PLD  devices) from  Altera.   Any
--other  use  of such  megafunction  design,  netlist,  support  information,
--device programming or simulation file,  or any other  related documentation
--or information  is prohibited  for  any  other purpose,  including, but not
--limited to  modification,  reverse engineering,  de-compiling, or use  with
--any other  silicon devices,  unless such use is  explicitly  licensed under
--a separate agreement with  Altera  or a megafunction partner.  Title to the
--intellectual property,  including patents,  copyrights,  trademarks,  trade
--secrets,  or maskworks,  embodied in any such megafunction design, netlist,
--support  information,  device programming or simulation file,  or any other
--related documentation or information provided by  Altera  or a megafunction
--partner, remains with Altera, the megafunction partner, or their respective
--licensors. No other licenses, including any licenses needed under any third
--party's intellectual property, are provided herein.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY cmd_queue_ram40 IS
	PORT
	(
		data		: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
		wraddress		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		rdaddress_a		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		rdaddress_b		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		wren		: IN STD_LOGIC  := '1';
		clock		: IN STD_LOGIC ;
		enable		: IN STD_LOGIC  := '1';
		qa		: OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
		qb		: OUT STD_LOGIC_VECTOR (39 DOWNTO 0)
	);
END cmd_queue_ram40;


ARCHITECTURE SYN OF cmd_queue_ram40 IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (39 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (39 DOWNTO 0);



	COMPONENT alt3pram
	GENERIC (
		intended_device_family		: STRING;
		width		: NATURAL;
		widthad		: NATURAL;
		indata_reg		: STRING;
		write_reg		: STRING;
		rdaddress_reg_a		: STRING;
		rdaddress_reg_b		: STRING;
		rdcontrol_reg_a		: STRING;
		rdcontrol_reg_b		: STRING;
		outdata_reg_a		: STRING;
		outdata_reg_b		: STRING;
		indata_aclr		: STRING;
		write_aclr		: STRING;
		rdaddress_aclr_a		: STRING;
		rdaddress_aclr_b		: STRING;
		rdcontrol_aclr_a		: STRING;
		rdcontrol_aclr_b		: STRING;
		outdata_aclr_a		: STRING;
		outdata_aclr_b		: STRING;
		lpm_type		: STRING;
		ram_block_type		: STRING;
		lpm_hint		: STRING
	);
	PORT (
			qa	: OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
			qb	: OUT STD_LOGIC_VECTOR (39 DOWNTO 0);
			inclocken	: IN STD_LOGIC ;
			wren	: IN STD_LOGIC ;
			inclock	: IN STD_LOGIC ;
			data	: IN STD_LOGIC_VECTOR (39 DOWNTO 0);
			rdaddress_a	: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			wraddress	: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			rdaddress_b	: IN STD_LOGIC_VECTOR (7 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	qa    <= sub_wire0(39 DOWNTO 0);
	qb    <= sub_wire1(39 DOWNTO 0);

	alt3pram_component : alt3pram
	GENERIC MAP (
		intended_device_family => "Stratix",
		width => 40,
		widthad => 8,
		indata_reg => "INCLOCK",
		write_reg => "INCLOCK",
		rdaddress_reg_a => "INCLOCK",
		rdaddress_reg_b => "INCLOCK",
		rdcontrol_reg_a => "UNREGISTERED",
		rdcontrol_reg_b => "UNREGISTERED",
		outdata_reg_a => "UNREGISTERED",
		outdata_reg_b => "UNREGISTERED",
		indata_aclr => "OFF",
		write_aclr => "OFF",
		rdaddress_aclr_a => "OFF",
		rdaddress_aclr_b => "OFF",
		rdcontrol_aclr_a => "OFF",
		rdcontrol_aclr_b => "OFF",
		outdata_aclr_a => "OFF",
		outdata_aclr_b => "OFF",
		lpm_type => "alt3pram",
		ram_block_type => "AUTO",
		lpm_hint => "USE_EAB=ON"
	)
	PORT MAP (
		inclocken => enable,
		wren => wren,
		inclock => clock,
		data => data,
		rdaddress_a => rdaddress_a,
		wraddress => wraddress,
		rdaddress_b => rdaddress_b,
		qa => sub_wire0,
		qb => sub_wire1
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: WidthData NUMERIC "40"
-- Retrieval info: PRIVATE: WidthAddr NUMERIC "8"
-- Retrieval info: PRIVATE: Clock NUMERIC "0"
-- Retrieval info: PRIVATE: rden_a NUMERIC "0"
-- Retrieval info: PRIVATE: rden_b NUMERIC "0"
-- Retrieval info: PRIVATE: REGdata NUMERIC "1"
-- Retrieval info: PRIVATE: REGwrite NUMERIC "1"
-- Retrieval info: PRIVATE: REGrdaddress_a NUMERIC "1"
-- Retrieval info: PRIVATE: REGrdaddress_b NUMERIC "1"
-- Retrieval info: PRIVATE: REGrren_a NUMERIC "0"
-- Retrieval info: PRIVATE: REGrren_b NUMERIC "0"
-- Retrieval info: PRIVATE: REGqa NUMERIC "0"
-- Retrieval info: PRIVATE: REGqb NUMERIC "0"
-- Retrieval info: PRIVATE: enable NUMERIC "1"
-- Retrieval info: PRIVATE: CLRdata NUMERIC "0"
-- Retrieval info: PRIVATE: CLRwrite NUMERIC "0"
-- Retrieval info: PRIVATE: CLRrdaddress_a NUMERIC "0"
-- Retrieval info: PRIVATE: CLRrdaddress_b NUMERIC "0"
-- Retrieval info: PRIVATE: CLRrren_a NUMERIC "0"
-- Retrieval info: PRIVATE: CLRrren_b NUMERIC "0"
-- Retrieval info: PRIVATE: CLRqa NUMERIC "0"
-- Retrieval info: PRIVATE: CLRqb NUMERIC "0"
-- Retrieval info: PRIVATE: BlankMemory NUMERIC "1"
-- Retrieval info: PRIVATE: MIFfilename STRING ""
-- Retrieval info: PRIVATE: UseLCs NUMERIC "0"
-- Retrieval info: PRIVATE: RAM_BLOCK_TYPE NUMERIC "0"
-- Retrieval info: PRIVATE: MAXIMUM_DEPTH NUMERIC "0"
-- Retrieval info: PRIVATE: INIT_FILE_LAYOUT STRING "PORT_A"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix"
-- Retrieval info: CONSTANT: WIDTH NUMERIC "40"
-- Retrieval info: CONSTANT: WIDTHAD NUMERIC "8"
-- Retrieval info: CONSTANT: INDATA_REG STRING "INCLOCK"
-- Retrieval info: CONSTANT: WRITE_REG STRING "INCLOCK"
-- Retrieval info: CONSTANT: RDADDRESS_REG_A STRING "INCLOCK"
-- Retrieval info: CONSTANT: RDADDRESS_REG_B STRING "INCLOCK"
-- Retrieval info: CONSTANT: RDCONTROL_REG_A STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: RDCONTROL_REG_B STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: OUTDATA_REG_A STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: OUTDATA_REG_B STRING "UNREGISTERED"
-- Retrieval info: CONSTANT: INDATA_ACLR STRING "OFF"
-- Retrieval info: CONSTANT: WRITE_ACLR STRING "OFF"
-- Retrieval info: CONSTANT: RDADDRESS_ACLR_A STRING "OFF"
-- Retrieval info: CONSTANT: RDADDRESS_ACLR_B STRING "OFF"
-- Retrieval info: CONSTANT: RDCONTROL_ACLR_A STRING "OFF"
-- Retrieval info: CONSTANT: RDCONTROL_ACLR_B STRING "OFF"
-- Retrieval info: CONSTANT: OUTDATA_ACLR_A STRING "OFF"
-- Retrieval info: CONSTANT: OUTDATA_ACLR_B STRING "OFF"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "alt3pram"
-- Retrieval info: CONSTANT: RAM_BLOCK_TYPE STRING "AUTO"
-- Retrieval info: CONSTANT: LPM_HINT STRING "USE_EAB=ON"
-- Retrieval info: USED_PORT: data 0 0 40 0 INPUT NODEFVAL data[39..0]
-- Retrieval info: USED_PORT: qa 0 0 40 0 OUTPUT NODEFVAL qa[39..0]
-- Retrieval info: USED_PORT: qb 0 0 40 0 OUTPUT NODEFVAL qb[39..0]
-- Retrieval info: USED_PORT: wraddress 0 0 8 0 INPUT NODEFVAL wraddress[7..0]
-- Retrieval info: USED_PORT: rdaddress_a 0 0 8 0 INPUT NODEFVAL rdaddress_a[7..0]
-- Retrieval info: USED_PORT: rdaddress_b 0 0 8 0 INPUT NODEFVAL rdaddress_b[7..0]
-- Retrieval info: USED_PORT: wren 0 0 0 0 INPUT VCC wren
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL clock
-- Retrieval info: USED_PORT: enable 0 0 0 0 INPUT VCC enable
-- Retrieval info: CONNECT: @data 0 0 40 0 data 0 0 40 0
-- Retrieval info: CONNECT: qa 0 0 40 0 @qa 0 0 40 0
-- Retrieval info: CONNECT: qb 0 0 40 0 @qb 0 0 40 0
-- Retrieval info: CONNECT: @wraddress 0 0 8 0 wraddress 0 0 8 0
-- Retrieval info: CONNECT: @rdaddress_a 0 0 8 0 rdaddress_a 0 0 8 0
-- Retrieval info: CONNECT: @rdaddress_b 0 0 8 0 rdaddress_b 0 0 8 0
-- Retrieval info: CONNECT: @wren 0 0 0 0 wren 0 0 0 0
-- Retrieval info: CONNECT: @inclock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @inclocken 0 0 0 0 enable 0 0 0 0
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
