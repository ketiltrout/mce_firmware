-- Copyright (c) 2003 SCUBA-2 Project
--                  All Rights Reserved
--
--  THIS IS UNPUBLISHED PROPRIETARY SOURCE CODE OF THE SCUBA-2 Project
--  The copyright notice above does not evidence any
--  actual or intended publication of such source code.
--
--  SOURCE CODE IS PROVIDED "AS IS". ALL EXPRESS OR IMPLIED CONDITIONS,
--  REPRESENTATIONS, AND WARRANTIES, INCLUDING ANY IMPLIED WARRANT OF
--  MERCHANTABILITY, SATISFACTORY QUALITY, FITNESS FOR A PARTICULAR
--  PURPOSE, OR NON-INFRINGEMENT, ARE DISCLAIMED, EXCEPT TO THE EXTENT
--  THAT SUCH DISCLAIMERS ARE HELD TO BE LEGALLY INVALID.
--
-- For the purposes of this code the SCUBA-2 Project consists of the
-- following organisations.
--
-- UKATC, Royal Observatory, Blackford Hill Edinburgh EH9 3HJ
-- UBC,   University of British Columbia, Physics & Astronomy Department,
--        Vancouver BC, V6T 1Z1
--
--
-- dispatch_reply_transmit.vhd
--
-- Project:	      SCUBA-2
-- Author:	       Ernie Lin
-- Organisation:  UBC
--
-- Description:
-- Implements the reply transmitter for the dispatch block.
--
-- Revision history:
-- 
-- $Log$
--
-----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library components;
use components.component_pack.all;

library work;
use work.async_pack.all;
use work.dispatch_pack.all;

entity dispatch_reply_transmit is
port(clk_i      : in std_logic;
     comm_clk_i : in std_logic;
     rst_i      : in std_logic;		
     
     lvds_tx_o : out std_logic;
     
     reply_rdy_i : in std_logic;
     reply_ack_o : out std_logic;  -- reply sent, clear to send next
     
     -- Command header words:
     header0_i : in std_logic_vector(PACKET_WORD_WIDTH-1 downto 0);
     header1_i : in std_logic_vector(PACKET_WORD_WIDTH-1 downto 0);
     header2_i : in std_logic_vector(PACKET_WORD_WIDTH-1 downto 0);  -- pass/fail word
     
     -- Buffer interface:
     buf_data_i : in std_logic_vector(BUF_DATA_WIDTH-1 downto 0);
     buf_addr_o : out std_logic_vector(BUF_ADDR_WIDTH-1 downto 0));
end dispatch_reply_transmit;

architecture rtl of dispatch_reply_transmit is

type transmitter_states is (IDLE_TX, CALC_CRC_START, WORD_TX_SETUP, WORD_TX_BUSY, CRC_TX_SETUP, CRC_TX_BUSY, TX_DONE);
signal tx_pres_state : transmitter_states;
signal tx_next_state : transmitter_states;

signal lvds_tx_data : std_logic_vector(PACKET_WORD_WIDTH-1 downto 0);
signal lvds_tx_rdy  : std_logic;
signal lvds_tx_busy : std_logic;

signal word_count_ena : std_logic;
signal word_count_clr : std_logic;
signal word_count     : integer;

signal reply_size    : std_logic_vector(DATA_SIZE_WIDTH-1 downto 0);
signal reply_size_ld : std_logic;

signal reply_num_words : integer;

-- signals used in CRC datapath:

type crc_states is (IDLE_CRC, INITIALIZE_CRC, CALCULATE_CRC, CRC_WORD_DONE, LOAD_NEXT_WORD, CRC_ALL_DONE);
signal crc_pres_state : crc_states;
signal crc_next_state : crc_states;

signal data_shreg_ena : std_logic;
signal data_shreg_ld  : std_logic;
signal crc_cur_bit    : std_logic;
signal crc_word_in    : std_logic_vector(PACKET_WORD_WIDTH-1 downto 0);
signal crc_word_out   : std_logic_vector(PACKET_WORD_WIDTH-1 downto 0);

signal crc_input_sel : std_logic_vector(1 downto 0);
signal tx_input_sel  : std_logic;

signal crc_bit_count_clr : std_logic;
signal crc_bit_count     : integer;

signal crc_ena   : std_logic;
signal crc_clr   : std_logic;
signal crc_done  : std_logic;
signal crc_checksum  : std_logic_vector(31 downto 0);

signal crc_num_bits : integer;

signal crc_word_rdy : std_logic;

signal crc_start : std_logic;
signal transmit_busy : std_logic;
signal transmit_done : std_logic;

begin

   ---------------------------------------------------------               
   -- Register for data size parameter
   ---------------------------------------------------------
   
   data_size_reg : reg
   generic map(WIDTH => DATA_SIZE_WIDTH)
   port map(clk_i => clk_i,
            rst_i => rst_i,
            ena_i => reply_size_ld,
            reg_i => header0_i(DATA_SIZE'range),
            reg_o => reply_size);
            
   -- number of bits to be processed by CRC is (# of data words + 2 header words + 1 pass/fail word) * 32
   crc_num_bits <= conv_integer((reply_size + 3) & "00000");
   
   -- number of words in packet (not including CRC) is (# of data words + 2 header words + 1 pass/fail word)
   reply_num_words <= conv_integer(reply_size + 3);
   
            
   ---------------------------------------------------------
   -- LVDS transmitter
   ---------------------------------------------------------

   reply_tx: lvds_tx
   port map(clk_i      => clk_i,
            comm_clk_i => comm_clk_i,
            rst_i      => rst_i,
            dat_i      => lvds_tx_data,
            rdy_i      => lvds_tx_rdy,
            busy_o     => lvds_tx_busy,
            lvds_o     => lvds_tx_o);
            
                                 
   ---------------------------------------------------------
   -- CRC calculation
   ---------------------------------------------------------

   crc_data_reg : shift_reg
      generic map(WIDTH => PACKET_WORD_WIDTH)
      port map(clk_i      => clk_i,
               rst_i      => rst_i,
               ena_i      => data_shreg_ena,
               load_i     => data_shreg_ld,
               clr_i      => '0',
               shr_i      => '1',
               serial_i   => crc_cur_bit, 
               serial_o   => crc_cur_bit,
               parallel_i => crc_word_in,
               parallel_o => crc_word_out);
                  
   crc_bit_counter : counter
      generic map(MAX         => PACKET_WORD_WIDTH,
                  WRAP_AROUND => '0')
      port map(clk_i   => clk_i,
               rst_i   => rst_i,
               ena_i   => '1',
               load_i  => crc_bit_count_clr,
               count_i => 0,
               count_o => crc_bit_count);

   crc_calc : crc
      generic map(POLY_WIDTH => 32)
      port map(clk_i      => clk_i,
               rst_i      => rst_i,
               clr_i      => crc_clr,
               ena_i      => crc_ena,
               data_i     => crc_cur_bit,
               num_bits_i => crc_num_bits,
               poly_i     => CRC32,
               done_o     => crc_done,
               valid_o    => open,
               checksum_o => crc_checksum);
               
   -- CRC control FSM
   crc_stateFF: process(clk_i, rst_i)
   begin
      if(rst_i = '1') then
         crc_pres_state <= IDLE_CRC;
      elsif(clk_i'event and clk_i = '1') then
         crc_pres_state <= crc_next_state;
      end if;
   end process crc_stateFF;
   
   crc_stateNS: process(crc_pres_state, crc_start, crc_bit_count, crc_done, transmit_busy, transmit_done)
   begin
      case crc_pres_state is
         when IDLE_CRC =>       if(crc_start = '1') then
                                   crc_next_state <= INITIALIZE_CRC;  
                                else
                                   crc_next_state <= IDLE_CRC;
                                end if;
                                   
         when INITIALIZE_CRC => crc_next_state <= CALCULATE_CRC;
                                
         when CALCULATE_CRC =>  if(crc_bit_count = PACKET_WORD_WIDTH-1) then
                                   crc_next_state <= CRC_WORD_DONE;
                                else
                                   crc_next_state <= CALCULATE_CRC;
                                end if;
                          
         when CRC_WORD_DONE =>  if(transmit_busy = '0') then              -- wait until previous word has been sent
                                   if(crc_done = '1') then
                                      crc_next_state <= CRC_ALL_DONE;
                                   else
                                      crc_next_state <= LOAD_NEXT_WORD;
                                   end if;
                                else
                                   crc_next_state <= CRC_WORD_DONE;
                                end if;
         
         when LOAD_NEXT_WORD => if(transmit_busy = '1') then
                                   crc_next_state <= CALCULATE_CRC;
                                else
                                   crc_next_state <= LOAD_NEXT_WORD;
                                end if;
         
         when CRC_ALL_DONE =>   if(transmit_done = '1') then
                                   crc_next_state <= IDLE_CRC;
                                else
                                   crc_next_state <= CRC_ALL_DONE;
                                end if;
                                         
         when others =>         crc_next_state <= IDLE_CRC;
      end case;
   end process crc_stateNS;
   
   crc_stateOut: process(crc_pres_state)
   begin 
      data_shreg_ena    <= '0';
      data_shreg_ld     <= '0';  
      crc_bit_count_clr <= '0';
      crc_ena           <= '0';
      crc_clr           <= '0';
      crc_word_rdy      <= '0';
      
      case crc_pres_state is
         when INITIALIZE_CRC => data_shreg_ena    <= '1';
                                data_shreg_ld     <= '1';
                                crc_bit_count_clr <= '1';
                                crc_ena           <= '1';
                                crc_clr           <= '1';
                           
         when CALCULATE_CRC =>  data_shreg_ena    <= '1';
                                crc_ena           <= '1';
         
         when CRC_WORD_DONE =>  crc_word_rdy      <= '1';
         
         when LOAD_NEXT_WORD => data_shreg_ena    <= '1';
                                data_shreg_ld     <= '1';
                                crc_bit_count_clr <= '1';
                                
         when others =>         null;
      end case;
   end process crc_stateOut;


   ---------------------------------------------------------               
   -- Counters for transmitted words
   ---------------------------------------------------------   
   
   word_counter : counter
   generic map(MAX => MAX_DATA_WORDS + 3)   -- there are 3 header words in addition to the data words
   port map(clk_i   => clk_i,
            rst_i   => rst_i,
            ena_i   => word_count_ena,
            load_i  => word_count_clr,
            count_i => 0,
            count_o => word_count);
            
   buf_addr_o <= conv_std_logic_vector(word_count - 3, BUF_ADDR_WIDTH);              -- data words start at word 3, header words are words 0-2.
   
   ---------------------------------------------------------               
   -- Multiplexors for inputs to CRC and LVDS blocks
   ---------------------------------------------------------
   
   with crc_input_sel select
      crc_word_in <= header0_i when "00",
                     header1_i when "01",
                     header2_i when "10",
                     buf_data_i when others;
   
   with tx_input_sel select
      lvds_tx_data <= crc_word_out when '0',
                      crc_checksum when others;
                      
      
   ---------------------------------------------------------
   -- Transmit controller FSM
   ---------------------------------------------------------
   tx_stateFF: process(clk_i, rst_i)
   begin
      if(rst_i = '1') then
         tx_pres_state <= IDLE_TX;
      elsif(clk_i'event and clk_i = '1') then
         tx_pres_state <= tx_next_state;
      end if;
   end process tx_stateFF;
   
   tx_stateNS: process(tx_pres_state, reply_rdy_i, crc_word_rdy, lvds_tx_busy, word_count)
   begin
      case tx_pres_state is
         when IDLE_TX =>        if(reply_rdy_i = '1') then
                                   tx_next_state <= CALC_CRC_START;
                                else
                                   tx_next_state <= IDLE_TX;
                                end if;
                          
         when CALC_CRC_START => if(crc_word_rdy = '1') then
                                   tx_next_state <= WORD_TX_SETUP;
                                else
                                   tx_next_state <= CALC_CRC_START;
                                end if;
         
         when WORD_TX_SETUP =>  tx_next_state <= WORD_TX_BUSY;
         
         when WORD_TX_BUSY =>   if(lvds_tx_busy = '0') then
                                   if(word_count = reply_num_words) then
                                      tx_next_state <= CRC_TX_SETUP;
                                   else
                                      tx_next_state <= WORD_TX_SETUP;
                                   end if;
                                else
                                   tx_next_state <= WORD_TX_BUSY;
                                end if;
 
         when CRC_TX_SETUP =>   tx_next_state <= CRC_TX_BUSY;
         
         when CRC_TX_BUSY =>    if(lvds_tx_busy = '0') then
                                   tx_next_state <= TX_DONE;
                                else
                                   tx_next_state <= CRC_TX_BUSY;
                                end if;
                          
         when TX_DONE =>        tx_next_state <= IDLE_TX;
      end case;
   end process tx_stateNS;
   
   tx_stateOut: process(tx_pres_state, word_count)
   begin
      case word_count is
         when 0 =>      crc_input_sel <= "00";
         when 1 =>      crc_input_sel <= "01";
         when 2 =>      crc_input_sel <= "10";
         when others => crc_input_sel <= "11";
      end case;
                                            
      -- default values:
      tx_input_sel   <= '0';
      reply_size_ld  <= '0';
      word_count_ena <= '0';
      word_count_clr <= '0';
      lvds_tx_rdy    <= '0';
      crc_start      <= '0';
      transmit_busy  <= '0';
      transmit_done  <= '0';
      reply_ack_o    <= '0';
      
      case tx_pres_state is
         when IDLE_TX =>                    reply_size_ld  <= '1';
                                            word_count_ena <= '1';
                                            word_count_clr <= '1';
                                
         when CALC_CRC_START =>             crc_start      <= '1';
         
         when WORD_TX_SETUP =>              tx_input_sel   <= '0';
                                            word_count_ena <= '1';
                                            lvds_tx_rdy    <= '1';
                                
         when WORD_TX_BUSY | CRC_TX_BUSY => transmit_busy  <= '1';

         when CRC_TX_SETUP =>               tx_input_sel   <= '1';
                                            lvds_tx_rdy    <= '1';
   
         when TX_DONE =>                    transmit_done  <= '1';
                                            reply_ack_o    <= '1';
      end case;
   end process tx_stateOut;
   
end rtl;