-- megafunction wizard: %LPM_MULT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: lpm_mult 

-- ============================================================
-- File Name: fsfb_corr_multiplier.vhd
-- Megafunction Name(s):
--          lpm_mult
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 4.1 Build 208 09/10/2004 SP 2 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2004 Altera Corporation
--Any  megafunction  design,  and related netlist (encrypted  or  decrypted),
--support information,  device programming or simulation file,  and any other
--associated  documentation or information  provided by  Altera  or a partner
--under  Altera's   Megafunction   Partnership   Program  may  be  used  only
--to program  PLD  devices (but not masked  PLD  devices) from  Altera.   Any
--other  use  of such  megafunction  design,  netlist,  support  information,
--device programming or simulation file,  or any other  related documentation
--or information  is prohibited  for  any  other purpose,  including, but not
--limited to  modification,  reverse engineering,  de-compiling, or use  with
--any other  silicon devices,  unless such use is  explicitly  licensed under
--a separate agreement with  Altera  or a megafunction partner.  Title to the
--intellectual property,  including patents,  copyrights,  trademarks,  trade
--secrets,  or maskworks,  embodied in any such megafunction design, netlist,
--support  information,  device programming or simulation file,  or any other
--related documentation or information provided by  Altera  or a megafunction
--partner, remains with Altera, the megafunction partner, or their respective
--licensors. No other licenses, including any licenses needed under any third
--party's intellectual property, are provided herein.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY fsfb_corr_multiplier IS
   PORT
   (
      dataa    : IN STD_LOGIC_VECTOR (31 DOWNTO 0); 
      datab    : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
      result      : OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
   );
END fsfb_corr_multiplier;


ARCHITECTURE SYN OF fsfb_corr_multiplier IS

   SIGNAL sub_wire0  : STD_LOGIC_VECTOR (63 DOWNTO 0);



   COMPONENT lpm_mult
   GENERIC (
      lpm_widtha     : NATURAL;
      lpm_widthb     : NATURAL;
      lpm_widthp     : NATURAL;
      lpm_widths     : NATURAL;
      lpm_type    : STRING;
      lpm_representation      : STRING;
      lpm_hint    : STRING
   );
   PORT (
         dataa : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
         datab : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
         result   : OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
   );
   END COMPONENT;

BEGIN
   result    <= sub_wire0(63 DOWNTO 0);

   lpm_mult_component : lpm_mult
   GENERIC MAP (
      lpm_widtha => 32,
      lpm_widthb => 32,
      lpm_widthp => 64,
      lpm_widths => 1,
      lpm_type => "LPM_MULT",
      lpm_representation => "SIGNED",
      lpm_hint => "DEDICATED_MULTIPLIER_CIRCUITRY=YES,MAXIMIZE_SPEED=5"
   )
   PORT MAP (
      dataa => dataa,
      datab => datab,
      result => sub_wire0
   );



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: WidthA NUMERIC "32"
-- Retrieval info: PRIVATE: WidthB NUMERIC "32"
-- Retrieval info: PRIVATE: WidthS NUMERIC "1"
-- Retrieval info: PRIVATE: WidthP NUMERIC "64"
-- Retrieval info: PRIVATE: OptionalSum NUMERIC "0"
-- Retrieval info: PRIVATE: AutoSizeResult NUMERIC "1"
-- Retrieval info: PRIVATE: B_isConstant NUMERIC "0"
-- Retrieval info: PRIVATE: SignedMult NUMERIC "1"
-- Retrieval info: PRIVATE: ConstantB NUMERIC "0"
-- Retrieval info: PRIVATE: ValidConstant NUMERIC "0"
-- Retrieval info: PRIVATE: Latency NUMERIC "0"
-- Retrieval info: PRIVATE: aclr NUMERIC "0"
-- Retrieval info: PRIVATE: clken NUMERIC "0"
-- Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "2"
-- Retrieval info: PRIVATE: optimize NUMERIC "1"
-- Retrieval info: CONSTANT: LPM_WIDTHA NUMERIC "32"
-- Retrieval info: CONSTANT: LPM_WIDTHB NUMERIC "32"
-- Retrieval info: CONSTANT: LPM_WIDTHP NUMERIC "64"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "1"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MULT"
-- Retrieval info: CONSTANT: LPM_REPRESENTATION STRING "SIGNED"
-- Retrieval info: CONSTANT: LPM_HINT STRING "DEDICATED_MULTIPLIER_CIRCUITRY=YES,MAXIMIZE_SPEED=5"
-- Retrieval info: USED_PORT: dataa 0 0 32 0 INPUT NODEFVAL dataa[31..0]
-- Retrieval info: USED_PORT: result 0 0 64 0 OUTPUT NODEFVAL result[63..0]
-- Retrieval info: USED_PORT: datab 0 0 32 0 INPUT NODEFVAL datab[31..0]
-- Retrieval info: CONNECT: @dataa 0 0 32 0 dataa 0 0 32 0
-- Retrieval info: CONNECT: result 0 0 64 0 @result 0 0 64 0
-- Retrieval info: CONNECT: @datab 0 0 32 0 datab 0 0 32 0
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL fsfb_corr_multiplier.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fsfb_corr_multiplier.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fsfb_corr_multiplier.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fsfb_corr_multiplier.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fsfb_corr_multiplier_inst.vhd FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fsfb_corr_multiplier_waveforms.html TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fsfb_corr_multiplier_wave*.jpg FALSE
