-- Copyright (c) 2003 SCUBA-2 Project
--                  All Rights Reserved
--
--  THIS IS UNPUBLISHED PROPRIETARY SOURCE CODE OF THE SCUBA-2 Project
--  The copyright notice above does not evidence any
--  actual or intended publication of such source code.
--
--  SOURCE CODE IS PROVIDED "AS IS". ALL EXPRESS OR IMPLIED CONDITIONS,
--  REPRESENTATIONS, AND WARRANTIES, INCLUDING ANY IMPLIED WARRANT OF
--  MERCHANTABILITY, SATISFACTORY QUALITY, FITNESS FOR A PARTICULAR
--  PURPOSE, OR NON-INFRINGEMENT, ARE DISCLAIMED, EXCEPT TO THE EXTENT
--  THAT SUCH DISCLAIMERS ARE HELD TO BE LEGALLY INVALID.
--
-- For the purposes of this code the SCUBA-2 Project consists of the
-- following organisations.
--
-- UKATC, Royal Observatory, Blackford Hill Edinburgh EH9 3HJ
-- UBC,   University of British Columbia, Physics & Astronomy Department,
--        Vancouver BC, V6T 1Z1
--
--
-- dip_switch_pack.vhd
--
-- Project:	      SCUBA-2
-- Author:	       Ernie Lin
-- Organisation:  UBC
--
-- Description:
-- Package file for dip switch module
--
-- Revision history:
-- 
-- $Log: dip_switch_pack.vhd,v $
-- Revision 1.2  2004/05/06 18:20:18  erniel
-- removed constant DIP_SWITCH_BITS
-- updated component declaration
--
--
-----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

library sys_param;
use sys_param.wishbone_pack.all;

package dip_switch_pack is
  
   component dip_switch    
      generic(WIDTH : in integer range 1 to 16 := 4);
      port(dip_switch_i : in std_logic_vector(WIDTH-1 downto 0);
     
           -- wishbone signals:
           clk_i  : in std_logic;
           rst_i  : in std_logic;
           addr_i : in std_logic_vector(WB_ADDR_WIDTH - 1 downto 0);
           dat_i  : in std_logic_vector(WB_DATA_WIDTH - 1 downto 0);
           dat_o  : out std_logic_vector(WB_DATA_WIDTH - 1 downto 0);
           tga_i  : in std_logic_vector(WB_TAG_ADDR_WIDTH - 1 downto 0);
           we_i   : in std_logic;
           stb_i  : in std_logic;
           cyc_i  : in std_logic;
           rty_o  : out std_logic;
           ack_o  : out std_logic);
   end component;

end dip_switch_pack;