-- Copyright (c) 2003 SCUBA-2 Project
--                  All Rights Reserved

--  THIS IS UNPUBLISHED PROPRIETARY SOURCE CODE OF THE SCUBA-2 Project
--  The copyright notice above does not evidence any
--  actual or intended publication of such source code.

--  SOURCE CODE IS PROVIDED "AS IS". ALL EXPRESS OR IMPLIED CONDITIONS,
--  REPRESENTATIONS, AND WARRANTIES, INCLUDING ANY IMPLIED WARRANT OF
--  MERCHANTABILITY, SATISFACTORY QUALITY, FITNESS FOR A PARTICULAR
--  PURPOSE, OR NON-INFRINGEMENT, ARE DISCLAIMED, EXCEPT TO THE EXTENT
--  THAT SUCH DISCLAIMERS ARE HELD TO BE LEGALLY INVALID.

-- For the purposes of this code the SCUBA-2 Project consists of the
-- following organisations.

-- UKATC, Royal Observatory, Blackford Hill Edinburgh EH9 3HJ
-- UBC,   University of British Columbia, Physics & Astronomy Department,
--        Vancouver BC, V6T 1Z1

-- 
--
-- <revision control keyword substitutions e.g. $Id: cmd_translator_simple_cmd_fsm.vhd,v 1.7 2004/05/06 18:16:43 jjacob Exp $>
--
-- Project:	      SCUBA-2
-- Author:	       Jonathan Jacob
--
-- Organisation:  UBC
--
-- Description:  This module is the fibre command translator. 
-- 
-- 
--
-- Revision history:
-- 
-- <date $Date: 2004/05/06 18:16:43 $>	-		<text>		- <initials $Author: jjacob $>
--
-- $Log$
--
-- 
-----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library components;
use components.component_pack.all;

library work;
use work.issue_reply_pack.all;

library sys_param;
use sys_param.wishbone_pack.all;
use sys_param.general_pack.all;


entity cmd_translator_simple_cmd_fsm is

--generic(cmd_translator_ADDR               : std_logic_vector(WB_ADDR_WIDTH-1 downto 0) := EEPROM_ADDR  );

port(

     -- global inputs

      rst_i        : in     std_logic;
      clk_i        : in     std_logic;

      -- inputs from cmd_translator top level      

      card_addr_i       : in std_logic_vector (CARD_ADDR_BUS_WIDTH-1 downto 0);  -- specifies which card the command is targetting
      parameter_id_i    : in std_logic_vector (PAR_ID_BUS_WIDTH-1 downto 0);     -- comes from reg_addr_i, indicates which device(s) the command is targetting
      data_size_i       : in std_logic_vector (DATA_SIZE_BUS_WIDTH-1 downto 0);  -- data_size_i, indicates number of 16-bit words of data
      data_i            : in std_logic_vector (DATA_BUS_WIDTH-1 downto 0);       -- data will be passed straight thru in 16-bit words
      data_clk_i        : in std_logic;							                         -- for clocking out the data
      
      -- other inputs
      sync_pulse_i    : in std_logic;
      cmd_start_i : in std_logic;
      cmd_stop_i  : in std_logic;
  
      -- outputs to the macro-instruction arbiter
      card_addr_o       : out std_logic_vector (CARD_ADDR_BUS_WIDTH-1 downto 0);  -- specifies which card the command is targetting
      parameter_id_o    : out std_logic_vector (PAR_ID_BUS_WIDTH-1 downto 0);     -- comes from reg_addr_i, indicates which device(s) the command is targetting
      data_size_o       : out std_logic_vector (DATA_SIZE_BUS_WIDTH-1 downto 0);  -- data_size_i, indicates number of 16-bit words of data
      data_o            : out std_logic_vector (DATA_BUS_WIDTH-1 downto 0);       -- data will be passed straight thru in 16-bit words
      data_clk_o        : out std_logic;							                          -- for clocking out the data
      macro_instr_rdy_o : out std_logic;                                          -- ='1' when the data is valid, else it's '0'
      
 
      -- input from the macro-instruction arbiter
      ack_i             : in std_logic                   -- acknowledgment from the micro-instr arbiter that it is ready and has grabbed the data

      -- outputs to the reply_translator block
      
      

   ); 
     
end cmd_translator_simple_cmd_fsm;


architecture rtl of cmd_translator_simple_cmd_fsm is


   type state is (IDLE, ISSUE_CMD);
   
   signal current_state, next_state : state;
   --signal word_count : integer;
   signal word_count     : std_logic_vector (DATA_SIZE_BUS_WIDTH-1 downto 0);
   signal zero_vector    : std_logic_vector (DATA_SIZE_BUS_WIDTH-2 downto 0);
   signal one            : std_logic;

begin

------------------------------------------------------------------------
--
-- state sequencer
--
------------------------------------------------------------------------

--   process(clk_i, rst_i)
--   begin
--      if rst_i = '1' then
--         current_state <= IDLE;
--      elsif clk_i'event and clk_i = '1' then
--         current_state <= next_state;
--      end if;
--   end process;

------------------------------------------------------------------------
--
-- assign next state
--
------------------------------------------------------------------------

--   process(current_state, cmd_start_i, word_count, data_size_i)
--   begin
--      case current_state is
--         when IDLE =>
--            if cmd_start_i = '1' then
--               next_state <= ISSUE_CMD;
--            else
--               next_state <= IDLE;
--            end if;
--            
--         when ISSUE_CMD =>
--            if word_count >= data_size_i then
--               next_state <= IDLE;--ISSUE_CMD_DONE;
--            else
--               next_state <= ISSUE_CMD;
--            end if;
--            
----         when ISSUE_CMD_DONE =>
----            next_state <= IDLE;
--            
--         when others =>
--            next_state <= IDLE;
--            
--      end case;
-- 
--   end process;
--

------------------------------------------------------------------------
--
-- assign outputs
--
------------------------------------------------------------------------

--   process(cmd_start_i, current_state, data_size_i, card_addr_i, parameter_id_i,
--           data_i, data_clk_i, word_count) -- maybe include word_count, but may cause delta-cycle issue
--   begin
--      case current_state is
--         when IDLE =>
--         
--            if cmd_start_i = '1' then
--            
--               card_addr_o        <= card_addr_i;
--               parameter_id_o     <= parameter_id_i;
--               data_size_o        <= data_size_i;
--               data_o             <= data_i;
--               data_clk_o         <= data_clk_i;
--               macro_instr_rdy_o  <= '1';
--            
--               --word_count         <= word_count + 1;
--
--            else
--
--               card_addr_o        <= (others => '0');
--               parameter_id_o     <= (others => '0');
--               data_size_o        <= (others => '0');
--               data_o             <= (others => '0');
--               data_clk_o         <= '0';
--               macro_instr_rdy_o  <= '0';
--            
--               --word_count         <= (others => '0');
--
--            end if;
--         
--         when ISSUE_CMD =>
--         
--            if word_count >= data_size_i then
--            
--               card_addr_o        <= (others => '0');
--               parameter_id_o     <= (others => '0');
--               data_size_o        <= (others => '0');
--               data_o             <= (others => '0');
--               data_clk_o         <= '0';
--               macro_instr_rdy_o  <= '0';
--            
--               --word_count         <= (others => '0');
--
--            else            
--               -- outputs to the macro-instruction arbiter
--               card_addr_o        <= card_addr_i;
--               parameter_id_o     <= parameter_id_i;
--               data_size_o        <= data_size_i;
--               data_o             <= data_i;
--               data_clk_o         <= data_clk_i;
--               macro_instr_rdy_o  <= '1';
--            
--               --word_count         <= word_count + 1;
--               
--            end if;
--         
--
--            
----         when ISSUE_CMD_DONE =>
--       
--      end case;
--   
--   end process;
--


------------------------------------------------------------------------
--
-- asynchronous state machine. Reacts immediately, no next-state clocking process
--
------------------------------------------------------------------------

   process(cmd_start_i, data_size_i, card_addr_i, parameter_id_i,
           data_i, data_clk_i, word_count) -- maybe include word_count, but may cause delta-cycle issue
   begin
      case current_state is
         when IDLE =>
         
            if cmd_start_i = '1' then
            
               card_addr_o        <= card_addr_i;
               parameter_id_o     <= parameter_id_i;
               data_size_o        <= data_size_i;
               data_o             <= data_i;
               data_clk_o         <= data_clk_i;
               macro_instr_rdy_o  <= '1';
            
               --word_count         <= word_count + 1;
               
               current_state <= ISSUE_CMD;

            else

               card_addr_o        <= (others => '0');
               parameter_id_o     <= (others => '0');
               data_size_o        <= (others => '0');
               data_o             <= (others => '0');
               data_clk_o         <= '0';
               macro_instr_rdy_o  <= '0';
            
               --word_count         <= (others => '0');
               current_state <= IDLE;

            end if;
         
         when ISSUE_CMD =>
         
            if word_count > data_size_i then
            
               card_addr_o        <= (others => '0');
               parameter_id_o     <= (others => '0');
               data_size_o        <= (others => '0');
               data_o             <= (others => '0');
               data_clk_o         <= '0';
               macro_instr_rdy_o  <= '0';
            
               --word_count         <= (others => '0');
               
               current_state <= IDLE;

            else            
               -- outputs to the macro-instruction arbiter
               card_addr_o        <= card_addr_i;
               parameter_id_o     <= parameter_id_i;
               data_size_o        <= data_size_i;
               data_o             <= data_i;
               data_clk_o         <= data_clk_i;
               macro_instr_rdy_o  <= '1';
            
               --word_count         <= word_count + 1;
               current_state <= ISSUE_CMD;
               
            end if;
         

            
--         when ISSUE_CMD_DONE =>
       
      end case;
   
   end process;
 
 
 
 

 
 
------------------------------------------------------------------------
--
-- word count
--
------------------------------------------------------------------------ 
-- write a counter based on data_clk
   process (current_state, data_clk_i)
   begin
      case current_state is
         when IDLE =>
            word_count <= (others => '0');
         when ISSUE_CMD =>
            if data_clk_i'event and data_clk_i='1' then
               word_count <= word_count + 1;
            end if;
         when others =>
            word_count <= (others => '0');
      end case;
   end process;
   
      
end rtl;