-- Copyright (c) 2003 SCUBA-2 Project
--                  All Rights Reserved

--  THIS IS UNPUBLISHED PROPRIETARY SOURCE CODE OF THE SCUBA-2 Project
--  The copyright notice above does not evidence any
--  actual or intended publication of such source code.

--  SOURCE CODE IS PROVIDED "AS IS". ALL EXPRESS OR IMPLIED CONDITIONS,
--  REPRESENTATIONS, AND WARRANTIES, INCLUDING ANY IMPLIED WARRANT OF
--  MERCHANTABILITY, SATISFACTORY QUALITY, FITNESS FOR A PARTICULAR
--  PURPOSE, OR NON-INFRINGEMENT, ARE DISCLAIMED, EXCEPT TO THE EXTENT
--  THAT SUCH DISCLAIMERS ARE HELD TO BE LEGALLY INVALID.

-- For the purposes of this code the SCUBA-2 Project consists of the
-- following organisations.

-- UKATC, Royal Observatory, Blackford Hill Edinburgh EH9 3HJ
-- UBC,   University of British Columbia, Physics & Astronomy Department,
--        Vancouver BC, V6T 1Z1

-- 
--
-- <revision control keyword substitutions e.g. $Id: issue_reply.vhd,v 1.31 2004/12/09 01:56:22 bburger Exp $>
--
-- Project:       SCUBA-2
-- Author:        Jonathan Jacob
--
-- Organisation:  UBC
--
-- Description:  This module is the top level for receiving fibre commands, translating them into
-- instructions, and issuing them over the bus backplane. 
-- 
--
-- Revision history:
-- 
-- <date $Date: 2004/12/09 01:56:22 $> -     <text>      - <initials $Author: bburger $>
--
-- $Log: issue_reply.vhd,v $
-- Revision 1.31  2004/12/09 01:56:22  bburger
-- Bryce:  updated the port map on the reply_translator to match the entity
--
-- Revision 1.30  2004/12/04 02:03:38  bburger
-- Bryce:  fixing some problems associated with integrating the reply_queue
--
-- Revision 1.29  2004/11/30 22:58:47  bburger
-- Bryce:  reply_queue integration
--
-- Revision 1.28  2004/11/25 11:04:30  dca
-- internal_cmd_i added to reply_translator instantiation
--
-----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library components;
use components.component_pack.all;

library work;
use work.issue_reply_pack.all;
use work.cmd_queue_pack.all;
use work.cmd_queue_ram40_pack.all;
use work.sync_gen_pack.all;
use work.fibre_rx_pack.all;
use work.fibre_tx_pack.all;
use work.reply_translator_pack.all;
use work.cmd_translator_pack.all;
use work.reply_queue_pack.all;

library sys_param;
use sys_param.command_pack.all;

entity issue_reply is
   port(
      -- for testing
      debug_o           : out std_logic_vector (31 downto 0);

      -- global signals
      rst_i             : in std_logic;
      clk_i             : in std_logic;
      comm_clk_i        : in std_logic;
      mem_clk_i         : in std_logic;
      
      -- inputs from the bus backplane
      lvds_reply_ac_a   : in std_logic;  
      lvds_reply_bc1_a  : in std_logic;
      lvds_reply_bc2_a  : in std_logic;
      lvds_reply_bc3_a  : in std_logic;
      lvds_reply_rc1_a  : in std_logic;
      lvds_reply_rc2_a  : in std_logic;
      lvds_reply_rc3_a  : in std_logic; 
      lvds_reply_rc4_a  : in std_logic;
      lvds_reply_cc_a   : in std_logic;
      
      -- inputs from the fibre receiver 
      fibre_clkr_i      : in std_logic;
      rx_data_i         : in std_logic_vector (7 DOWNTO 0);
      nRx_rdy_i         : in std_logic;
      rvs_i             : in std_logic;
      rso_i             : in std_logic;
      rsc_nRd_i         : in std_logic;        
      cksum_err_o       : out std_logic;

      -- interface to fibre transmitter
      tx_data_o         : out std_logic_vector (7 downto 0);      -- byte of data to be transmitted
      tsc_nTd_o         : out std_logic;                          -- hotlink tx special char/ data sel
      nFena_o           : out std_logic;                           -- hotlink tx enable

      -- 25MHz clock for fibre_tx_control
      fibre_clkw_i      : in std_logic;                          -- in phase with 25MHz hotlink clock

      -- lvds_tx interface
      lvds_cmd_o              : out std_logic;  -- transmitter output pin

      -- sync_gen interface
      sync_pulse_i      : in std_logic;
      sync_number_i     : in std_logic_vector (SYNC_NUM_WIDTH-1 downto 0)
   );     
end issue_reply;


architecture rtl of issue_reply is

   -- inputs from fibre_rx 
   signal card_id             : std_logic_vector (FIBRE_CARD_ADDRESS_WIDTH-1 downto 0);    -- specifies which card the command is targetting
   signal cmd_code            : std_logic_vector (15 downto 0);                       -- the least significant 16-bits from the fibre packet
   signal cksum_err           : std_logic;
   signal cmd_data            : std_logic_vector (PACKET_WORD_WIDTH-1 downto 0);         -- the data 
   signal cmd_rdy             : std_logic;                                            -- indicates the fibre_rx outputs are valid
   signal data_clk            : std_logic;                                            -- used to clock the data out
   signal num_data            : std_logic_vector (FIBRE_DATA_SIZE_WIDTH-1 downto 0);    -- number of 16-bit data words to be clocked out, possibly number of bytes
   signal param_id            : std_logic_vector (FIBRE_PARAMETER_ID_WIDTH-1 downto 0);       -- the parameter ID
   signal cmd_type            : std_logic_vector (BB_COMMAND_TYPE_WIDTH-1 downto 0);       -- this is a re-mapping of the cmd_code into a 3-bit number
   signal cmd_ack             : std_logic;   -- acknowledge signal from cmd_translator to fibre_rx
  
   signal reply_cmd_rcvd_er   : std_logic;
   signal reply_cmd_rcvd_ok   : std_logic;
   signal reply_cmd_code      : std_logic_vector (15 downto 0);
   signal reply_param_id      : std_logic_vector (FIBRE_PARAMETER_ID_WIDTH-1 downto 0); 
   signal reply_card_id       : std_logic_vector (FIBRE_CARD_ADDRESS_WIDTH-1 downto 0);

   signal sync_pulse          : std_logic;
   signal sync_number         : std_logic_vector (7 downto 0);
   
   -- reply_queue interface
   signal uop_status          : std_logic_vector(BB_STATUS_WIDTH-1 downto 0);
   signal uop_rdy             : std_logic;
   signal uop_rdy_stg1        : std_logic;
   signal uop_rdy_stg2        : std_logic;
   signal uop_rdy_stg3        : std_logic;
   signal uop_rdy_stg4        : std_logic;
   signal uop_rdy_stg5        : std_logic;
   
   signal uop_ack             : std_logic;
   signal uop_discard         : std_logic;
   signal uop_timedout        : std_logic;
   signal uop                 : std_logic_vector(QUEUE_WIDTH-1 downto 0);  
 
   -- cmd_translator to cmd_queue interface
   signal card_addr           : std_logic_vector (FIBRE_CARD_ADDRESS_WIDTH-1 downto 0);
   signal parameter_id        : std_logic_vector (FIBRE_PARAMETER_ID_WIDTH-1 downto 0); 
   signal data_size           : std_logic_vector (FIBRE_DATA_SIZE_WIDTH-1 downto 0);
   signal data                : std_logic_vector (PACKET_WORD_WIDTH-1 downto 0);
   signal data_clk2           : std_logic; 
   signal m_op_seq_num        : std_logic_vector(BB_MACRO_OP_SEQ_WIDTH-1 downto 0);
   signal frame_sync_num      : std_logic_vector(SYNC_NUM_WIDTH-1 downto 0);
   signal frame_seq_num       : std_logic_vector(PACKET_WORD_WIDTH-1 downto 0);
   signal macro_instr_rdy     : std_logic; 
   signal mop_ack             : std_logic; 
   signal cmd_stop            : std_logic;
   signal last_frame          : std_logic;      
   signal internal_cmd_issued : std_logic;
   
   -- reply_translator to reply_queue interface      
   signal m_op_rdy            : std_logic;     
   signal m_op_error_code     : std_logic_vector(29 downto 0); 
   signal m_op_cmd_code       : std_logic_vector(BB_COMMAND_TYPE_WIDTH-1    downto 0); 
   signal m_op_param_id       : std_logic_vector (BB_PARAMETER_ID_WIDTH-1  downto 0);  
   signal m_op_card_id        : std_logic_vector (BB_CARD_ADDRESS_WIDTH-1  downto 0);  
   signal fibre_word          : std_logic_vector (PACKET_WORD_WIDTH-1        downto 0); 
   signal num_fibre_words     : integer;    
   signal fibre_word_ack      : std_logic;
   signal fibre_word_rdy      : std_logic;
   signal m_op_ack            : std_logic;   
   signal reply_cmd_stop      : std_logic;
   signal reply_last_frame    : std_logic;
   signal reply_frame_seq_num : std_logic_vector(PACKET_WORD_WIDTH-1 downto 0);
   signal internal_cmd        : std_logic := '0';
 
   -- reply_translator / fibre_tx interface 
   signal txd                 : std_logic_vector(7 downto 0); 
   signal tx_fw               : std_logic; 
   signal tx_ff               : std_logic;     
   
   type state is (IDLE, WAIT1, WAIT2, ACK1, ACK2);
   signal cur_state, next_state  : state;

begin
   -- temporarily routing these signals to top level to view them on the logic analyzer
--   parameter_id_o    <= parameter_id;
--   data_o            <= data;
--   data_clk_o        <= data_clk2;
--   macro_instr_rdy_o <= cmd_rdy;
--   macro_op_ack_o    <= cmd_ack;

   ------------------------------------------------------------------------
   -- fibre receiver
   ------------------------------------------------------------------------
   i_fibre_rx : fibre_rx
      port map( 
         rst_i        => rst_i,
         clk_i        => clk_i,
         
         -- inputs from the fibre
         fibre_clkr_i => fibre_clkr_i,
         nrx_rdy_i    => nrx_rdy_i,
         rvs_i        => rvs_i,
         rso_i        => rso_i,
         rsc_nrd_i    => rsc_nrd_i,
         rx_data_i    => rx_data_i,
         
         -- input from cmd_translator
         cmd_ack_i    => cmd_ack,                  -- command acknowledge
         
         -- outputs to cmd_translator
         cmd_code_o   => cmd_code,                   -- command code
         card_id_o    => card_id,                    -- card id
         param_id_o   => param_id,                   -- parameter id
         num_data_o   => num_data,                   -- number of valid 32 bit data words
         cmd_data_o   => cmd_data,                   -- 32bit valid data word
         cmd_rdy_o    => cmd_rdy,                    -- checksum error flag
         data_clk_o   => data_clk,                   -- data clock
         
         cksum_err_o  => cksum_err
      );

   cksum_err_o <= cksum_err;

   ------------------------------------------------------------------------
   -- fibre transmitter
   ------------------------------------------------------------------------
   i_fibre_tx : fibre_tx
      port map(        
         -- global inputs
         clk_i        => clk_i, 
         rst_i        => rst_i, 
            
         -- interface to reply_translator 
         txd_i        => txd, 
         tx_fw_i      => tx_fw, 
         tx_ff_o      => tx_ff, 
         
         -- interface to HOTLINK transmitter
         fibre_clkw_i => fibre_clkw_i,
         tx_data_o    => tx_data_o,
         tsc_nTd_o    => tsc_nTd_o,
         nFena_o      => nFena_o 
      );

   ------------------------------------------------------------------------
   -- reply_translator
   ------------------------------------------------------------------------ 
   i_reply_translator : reply_translator
      port map(
         -- global inputs 
         rst_i             => rst_i,
         clk_i             => clk_i,

         -- signals to/from cmd_translator    
         cmd_rcvd_er_i     => reply_cmd_rcvd_er,
         cmd_rcvd_ok_i     => reply_cmd_rcvd_ok,
         cmd_code_i        => reply_cmd_code,
         card_id_i         => reply_card_id,
         param_id_i        => reply_param_id,            
                         
         -- signals to/from reply queue
         mop_rdy_i        => m_op_rdy,  
         mop_error_code_i => m_op_error_code, 
         mop_cmd_code_i   => m_op_cmd_code,
         mop_param_id_i   => m_op_param_id,
         mop_card_id_i    => m_op_card_id, 
         internal_cmd_i    => internal_cmd,
         fibre_word_i      => fibre_word,
         num_fibre_words_i => num_fibre_words,
         fibre_word_ack_o  => fibre_word_ack,
         fibre_word_rdy_i  => fibre_word_rdy,
         mop_ack_o        => m_op_ack,    
         
         cmd_stop_i        => reply_cmd_stop,
         last_frame_i      => reply_last_frame,
         frame_seq_num_i   => reply_frame_seq_num,

         -- signals to / from fibre_tx
         tx_ff_i           => tx_ff, 
         tx_fw_o           => tx_fw,
         txd_o             => txd
      );      

   ------------------------------------------------------------------------
   -- command translator
   ------------------------------------------------------------------------
   i_cmd_translator : cmd_translator
      port map(
         -- global inputs
         rst_i               => rst_i,
         clk_i               => clk_i,
         
         -- inputs from fibre_rx
         card_id_i           => card_id,
         cmd_code_i          => cmd_code,
         cmd_data_i          => cmd_data,
         cksum_err_i         => cksum_err,
         cmd_rdy_i           => cmd_rdy,
         data_clk_i          => data_clk,
         num_data_i          => num_data,
         param_id_i          => param_id,
         
         -- output to fibre_rx
         ack_o               => cmd_ack,
         
         -- outputs to u-op sequence generator         
         card_addr_o         => card_addr,--card_addr_o,
         parameter_id_o      => parameter_id,--parameter_id_o,
         data_size_o         => data_size,--data_size_o,
         data_o              => data,--data_o,
         data_clk_o          => data_clk2,--data_clk_o,
         macro_instr_rdy_o   => macro_instr_rdy,--macro_instr_rdy_o,
         m_op_seq_num_o      => m_op_seq_num,--m_op_seq_num_o,
         frame_seq_num_o     => frame_seq_num,--frame_seq_num_o,
         frame_sync_num_o    => frame_sync_num,--frame_sync_num_o,
         cmd_type_o          => cmd_type,
         cmd_stop_o          => cmd_stop,
         last_frame_o        => last_frame,       
         internal_cmd_o      => internal_cmd_issued,
         
         --input from the u-op sequence generator
         ack_i               => mop_ack,
         
         -- reply_translator interface          
         reply_cmd_rcvd_er_o => reply_cmd_rcvd_er,
         reply_cmd_rcvd_ok_o => reply_cmd_rcvd_ok,
         reply_cmd_code_o    => reply_cmd_code,
         reply_param_id_o    => reply_param_id,
         reply_card_id_o     => reply_card_id,         
         
         sync_pulse_i        => sync_pulse_i,
         sync_number_i       => sync_number_i
      );

   ------------------------------------------------------------------------
   -- command queue (u-op sequence generator)
   ------------------------------------------------------------------------               
   uop_status <= (others=>'0');
     
   i_cmd_queue : cmd_queue
     port map(
        -- for testing
        debug_o         => debug_o,

        -- reply_queue interface
        uop_rdy_o       => uop_rdy,
        uop_ack_i       => uop_ack,  --uop_rdy_stg5
        uop_o           => uop,
        
        -- cmd_translator interface
        card_addr_i     => card_addr,
        par_id_i        => parameter_id,
        data_size_i     => data_size,
        data_i          => data,
        data_clk_i      => data_clk2,
        mop_i           => m_op_seq_num,
        issue_sync_i    => frame_sync_num,
        mop_rdy_i       => macro_instr_rdy,
        mop_ack_o       => mop_ack,
        cmd_type_i      => cmd_type,
        cmd_stop_i      => cmd_stop,
        last_frame_i    => last_frame,
        frame_seq_num_i => frame_seq_num,--frame_seq_num_o,
        internal_cmd_i  => internal_cmd_issued,

        -- lvds_tx interface
        tx_o            => lvds_cmd_o,

        -- frame_timing interface
        sync_i          => sync_pulse_i,
        sync_num_i      => sync_number_i,

        -- Clock lines
        clk_i           => clk_i,
        comm_clk_i      => comm_clk_i,
        mem_clk_i       => mem_clk_i,
        rst_i           => rst_i
     );

   ------------------------------------------------------------------------
   -- reply queue
   ------------------------------------------------------------------------
   i_reply_queue : reply_queue
      port map(
         -- cmd_queue interface
         cmd_to_retire_i  => uop_rdy,
         cmd_sent_o       => uop_ack,
         cmd_i            => uop,
         
         -- reply_translator interface (from reply_queue, i.e. these signals are de-multiplexed from retire and sequencer)
         size_o           => num_fibre_words,
         data_o           => fibre_word,
         error_code_o     => m_op_error_code,
         cmd_valid_o      => m_op_rdy,
         rdy_o            => fibre_word_rdy,
         ack_i            => fibre_word_ack,
         
         -- reply_translator interface (from reply_queue_retire)
         cmd_sent_i       => m_op_ack,
         cmd_code_o       => m_op_cmd_code,
         param_id_o       => m_op_param_id,
         card_addr_o      => m_op_card_id,
         stop_bit_o       => reply_cmd_stop,
         last_frame_bit_o => reply_last_frame,
         frame_seq_num_o  => reply_frame_seq_num,
         internal_cmd_o   => internal_cmd,
   
         -- Bus Backplane interface
         lvds_reply_ac_a     => lvds_reply_ac_a,
         lvds_reply_bc1_a    => lvds_reply_bc1_a,
         lvds_reply_bc2_a    => lvds_reply_bc2_a,
         lvds_reply_bc3_a    => lvds_reply_bc3_a,
         lvds_reply_rc1_a    => lvds_reply_rc1_a,
         lvds_reply_rc2_a    => lvds_reply_rc2_a,
         lvds_reply_rc3_a    => lvds_reply_rc3_a,
         lvds_reply_rc4_a    => lvds_reply_rc4_a,
         lvds_reply_cc_a     => lvds_reply_cc_a,
         
         -- Global signals
         clk_i            => clk_i,
         mem_clk_i        => mem_clk_i,
         comm_clk_i       => comm_clk_i,
         rst_i            => rst_i
      );

end rtl; 