-- Copyright (c) 2003 SCUBA-2 Project
-- All Rights Reserved
-- THIS IS UNPUBLISHED PROPRIETARY SOURCE CODE OF THE SCUBA-2 Project
-- The copyright notice above does not evidence any
-- actual or intended publication of such source code.
-- SOURCE CODE IS PROVIDED "AS IS". ALL EXPRESS OR IMPLIED CONDITIONS,
-- REPRESENTATIONS, AND WARRANTIES, INCLUDING ANY IMPLIED WARRANT OF
-- MERCHANTABILITY, SATISFACTORY QUALITY, FITNESS FOR A PARTICULAR
-- PURPOSE, OR NON-INFRINGEMENT, ARE DISCLAIMED, EXCEPT TO THE EXTENT
-- THAT SUCH DISCLAIMERS ARE HELD TO BE LEGALLY INVALID.
-- For the purposes of this code the SCUBA-2 Project consists of the
-- following organisations.
-- UKATC, Royal Observatory, Blackford Hill Edinburgh EH9 3HJ
-- UBC, University of British Columbia, Physics & Astronomy Department,
-- Vancouver BC, V6T 1Z1
-- 
--
--
-- Project:      Scuba 2
-- Author:       Mandana Amiri
-- Organisation: UBC
-- original source: tb_bias_card_self_test
-- revised by:   Mandana Amiri
--
-- Title
-- tb_bias_card_self_test
--
-- Description:
-- Revision history:
-- <date $Date: 2006/03/02 19:05:06 $>    - <initials $Author: mandana $>
-- $Log: tb_bias_card_self_test.vhd,v $
-- Revision 1.4  2006/03/02 19:05:06  mandana
-- took out non-bias-card related signals
--
-- Revision 1.3  2005/02/01 01:09:39  mandana
-- slot_id and ttl_nrx1 are now hard coded in the self_test module
--
-- Revision 1.2  2005/01/27 00:13:38  mandana
-- ttl_nrx, ttl_tx, ttl_txena changed from vector to std_logic!
--
-- Revision 1.1  2005/01/20 22:49:14  mandana
-- Inital Release: bias_card self-test with incoming packets pushed in from the RAM
--   
--
-------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

library work;
use work.bc_dac_ctrl_pack.all;
use work.clk_card_pack.all;
use work.bias_card_pack.all;
use work.addr_card_pack.all;

library components;
use components.component_pack.all;

library sys_param;
use sys_param.command_pack.all;
use sys_param.wishbone_pack.all;
use sys_param.data_types_pack.all;

entity tb_bias_card_self_test is     
end tb_bias_card_self_test;

architecture tb of tb_bias_card_self_test is 
 

   constant clk_period     : TIME := 40 ns;    -- 25Mhz clock input to PLL
   constant clk_spi_period : TIME := 40 ns;    -- 25MHz clock
        
   constant flux_fdbck_cmd : std_logic_vector(31 downto 0) := x"00" & BIAS_CARD_1        & x"00" & FLUX_FB_ADDR;
   constant bias_cmd       : std_logic_vector(31 downto 0) := x"00" & BIAS_CARD_1        & x"00" & BIAS_ADDR;
   constant led_cmd        : std_logic_vector(31 downto 0) := x"00" & BIAS_CARD_1        & x"00" & LED_ADDR;
   constant sram1_strt_cmd : std_logic_vector(31 downto 0) := x"00" & CLOCK_CARD         & x"00" & SRAM1_STRT_ADDR;  
         
   ------------------------------------------------
   -- Bias Card Signals
   -------------------------------------------------    
   signal   rst_n       : std_logic := '1';   
   signal   inclk       : std_logic := '0';
   
   -- lvds signals
   signal lvds_sync     : std_logic := '0'; --52us clock, normally generated by clock_card/sync_gen block, but testbench generated here
   signal lvds_spare    : std_logic;
   signal lvds_reply_bc1_a : std_logic := '0';
   signal lvds_reply_bc1_b : std_logic := '0';
   
   -- TTL interface:
   signal ttl_nrx1      : std_logic;
   signal ttl_tx1       : std_logic;
   signal ttl_txena1    : std_logic;
		       
   signal ttl_nrx2      : std_logic;
   signal ttl_tx2       : std_logic;
   signal ttl_txena2    : std_logic;
		       
   signal ttl_nrx3      : std_logic;
   signal ttl_tx3       : std_logic;
   signal ttl_txena3    : std_logic;
   		       
   -- eeprom interface:
   signal bc_eeprom_si  : std_logic := '0';
   signal bc_eeprom_so  : std_logic;
   signal bc_eeprom_sck : std_logic;
   signal bc_eeprom_cs  : std_logic;
    
   -- dac interface:
   signal dac_ncs       : std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);
   signal dac_sclk      : std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);
   signal dac_data      : std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);      
   signal lvds_dac_ncs  : std_logic;
   signal lvds_dac_sclk : std_logic;
   signal lvds_dac_data : std_logic;
   signal dac_nclr      : std_logic; -- add to tcl file
   
   -- miscellaneous ports:
   signal bc_red_led    : std_logic;
   signal bc_ylw_led    : std_logic;
   signal bc_grn_led    : std_logic;
   signal bc_dip_sw3    : std_logic;
   signal bc_dip_sw4    : std_logic;
   signal bc_wdog       : std_logic;
   signal bc_slot_id    : std_logic_vector(3 downto 0) := "1110";
    
   -- debug ports:
   signal bc_rs232_rx   : std_logic;
   signal bc_rs232_tx   : std_logic;   
   signal test          : std_logic_vector(16 downto 3);
   signal mictor        : std_logic_vector(32 downto 1);
   signal mictorclk     : std_logic_vector(2 downto 1);
   		        
   -- simulation signals
   signal pdat          : std_logic_vector(7 downto 0) := x"00";   
   
   -- RAM containing the backplane instructions
   component packet_ram
   	PORT
   	(
   		address		: IN STD_LOGIC_VECTOR (5 DOWNTO 0);
   		clock		: IN STD_LOGIC ;
   		data		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
   		wren		: IN STD_LOGIC ;
   		q		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
   	);
   end component;
   
begin
  
   i_bias_card_self_test: bias_card_self_test
      port map(

         -- PLL input:
         inclk      => inclk,
         rst_n      => rst_n,
         
         -- LVDS interface:
 --        lvds_cmd   => lvds_lvds_tx, --lvds_cmd,  
         lvds_sync  => lvds_sync, 
         lvds_spare => lvds_spare,
         lvds_txa   => lvds_reply_bc1_a, 
         lvds_txb   => lvds_reply_bc1_b, 
         
         -- TTL interface:
--        ttl_nrx1    => ttl_nrx1,  
         ttl_tx1     => ttl_tx1,   
         ttl_txena1  => ttl_txena1,

         ttl_nrx2    => ttl_nrx2,  
         ttl_tx2     => ttl_tx2,   
         ttl_txena2  => ttl_txena2,

         ttl_nrx3    => ttl_nrx3,  
         ttl_tx3     => ttl_tx3,   
         ttl_txena3  => ttl_txena3,
         
         -- eeprom ice:nterface:
         eeprom_si  => bc_eeprom_si, 
         eeprom_so  => bc_eeprom_so, 
         eeprom_sck => bc_eeprom_sck,
         eeprom_cs  => bc_eeprom_cs, 
         
         -- dac interface:
         dac_ncs    => dac_ncs,      
         dac_sclk   => dac_sclk,     
         dac_data   => dac_data,         
         lvds_dac_ncs  => lvds_dac_ncs, 
         lvds_dac_sclk => lvds_dac_sclk,
         lvds_dac_data => lvds_dac_data,
         dac_nclr      => dac_nclr,     
         
         -- miscellaneous ports:
         red_led    => bc_red_led, 
         ylw_led    => bc_ylw_led, 
         grn_led    => bc_grn_led, 
         dip_sw3    => bc_dip_sw3, 
         dip_sw4    => bc_dip_sw4, 
         wdog       => bc_wdog,    
--         slot_id    => bc_slot_id, 
         
         -- debug ports:
         test       => test,       
         mictor     => mictor,     
         mictorclk  => mictorclk,  
         rx   => bc_rs232_rx,
         tx   => bc_rs232_tx
      );     
      
    --   bc_slot_id      <= "1110";
    --   cc_slot_id      <= "1000";
   ------------------------------------------------
   -- Create test bench clock
   -------------------------------------------------
   --   ttl_nrx1     <= '0';
   inclk        <= not inclk        after clk_period/2;   
   lvds_sync    <= not lvds_sync    after clk_period*2600/2;   
   
   ------------------------------------------------------------------------------
   -- emulate external interface
   --
   emulate_ee_data: process -- emulate data read from eeprom on the spi_si line
   begin
      wait until bc_eeprom_cs = '0';
      wait for 33*clk_period;
      for j in 0 to 5 loop
         pdat <= pdat + 23;
         wait for 6*clk_period;
         for i in 0 to 7 loop      
           bc_eeprom_si <= pdat(7-i);  
           wait for clk_spi_period;      
         end loop;
      end loop;
   end process emulate_ee_data;   

   ------------------------------------------------
   -- Create test bench stimuli
   -------------------------------------------------
   stimuli : process
   procedure do_reset is
   begin
      rst_n <= '0';
      wait for clk_period*5 ;
      rst_n <= '1';
      wait for clk_period*5 ;   
      assert false report " Resetting the DUT." severity NOTE;
   end do_reset;
  
--------------------------------------------------------
-- Begin Test
------------------------------------------------------      
   begin
      
      do_reset;                
      wait for 120 us;
      assert false report "Simulation done." severity FAILURE;
   end process stimuli;   
end tb;