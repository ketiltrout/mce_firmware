-- 2003 SCUBA-2 Project
--                  All Rights Reserved

--  THIS IS UNPUBLISHED PROPRIETARY SOURCE CODE OF THE SCUBA-2 Project
--  The copyright notice above does not evidence any
--  actual or intended publication of such source code.

--  SOURCE CODE IS PROVIDED "AS IS". ALL EXPRESS OR IMPLIED CONDITIONS,
--  REPRESENTATIONS, AND WARRANTIES, INCLUDING ANY IMPLIED WARRANT OF
--  MERCHANTABILITY, SATISFACTORY QUALITY, FITNESS FOR A PARTICULAR
--  PURPOSE, OR NON-INFRINGEMENT, ARE DISCLAIMED, EXCEPT TO THE EXTENT
--  THAT SUCH DISCLAIMERS ARE HELD TO BE LEGALLY INVALID.

-- For the purposes of this code the SCUBA-2 Project consists of the
-- following organisations.

-- UKATC, Royal Observatory, Blackford Hill Edinburgh EH9 3HJ
-- UBC,   University of British Columbia, Physics & Astronomy Department,
--        Vancouver BC, V6T 1Z1

-- $Id: bc_dac_ctrl.vhd,v 1.7 2006/08/03 19:06:31 mandana Exp $
--
-- Project:       SCUBA2
-- Author:        Bryce Burger
-- Organisation:  UBC
--
-- Description:
-- This block processes wishbone commands FLUX_FB_ADDR and BIAS_ADDR and 
-- updates 32 flux_fb SPI DACs and 12 low-noise bias SPI DACs.
-- 
-- Revision history:
-- $Log: bc_dac_ctrl.vhd,v $
-- Revision 1.7  2006/08/03 19:06:31  mandana
-- reorganized pack files, bc_dac_ctrl_core_pack, bc_dac_ctrl_wbs_pack, frame_timing_pack are all obsolete
--
-- Revision 1.6  2005/01/17 23:01:04  mandana
-- removed mem_clk_i
-- read from RAM is performed in 2 clk_i cycles, added an extra state for read
--
-- Revision 1.5  2005/01/04 19:19:47  bburger
-- Mandana: changed mictor assignment to 0 to 31 and swapped odd and even pods
--
-- Revision 1.4  2004/12/21 22:06:51  bburger
-- Bryce:  update
--
-- Revision 1.3  2004/11/25 03:05:08  bburger
-- Bryce:  Modified the Bias Card DAC control slaves.
--
-- Revision 1.2  2004/11/15 20:03:41  bburger
-- Bryce :  Moved frame_timing to the 'work' library, and physically moved the files to "all_cards" directory
--
-- Revision 1.1  2004/11/11 01:47:10  bburger
-- Bryce:  new
--
--   
--
-- 
-----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

library sys_param;
use sys_param.wishbone_pack.all;

library work;
use work.bias_card_pack.all;
use work.bc_dac_ctrl_pack.all;

entity bc_dac_ctrl is
   port
   (
      -- DAC hardware interface:
      -- 32 independant flux-fb DAC channels, thus 32 serial data/cs/clk lines and
      -- 12 ln_bias DAC channels, data and clk lines are shared
      flux_fb_data_o    : out std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);   
      flux_fb_ncs_o     : out std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);
      flux_fb_clk_o     : out std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);      
      
      ln_bias_data_o    : out std_logic;
      ln_bias_ncs_o     : out std_logic_vector(NUM_LN_BIAS_DACS-1 downto 0);
      ln_bias_clk_o     : out std_logic;
      
      dac_nclr_o        : out std_logic;
      
      -- wishbone interface:
      dat_i             : in std_logic_vector(WB_DATA_WIDTH-1 downto 0);
      addr_i            : in std_logic_vector(WB_ADDR_WIDTH-1 downto 0);
      tga_i             : in std_logic_vector(WB_TAG_ADDR_WIDTH-1 downto 0);
      we_i              : in std_logic;
      stb_i             : in std_logic;
      cyc_i             : in std_logic;
      dat_o             : out std_logic_vector(WB_DATA_WIDTH-1 downto 0);
      ack_o             : out std_logic;
      
      -- frame_timing signals
      update_bias_i     : in std_logic;
      restart_frame_aligned_i : in std_logic;      
      
      -- Global Signals      
      clk_i             : in std_logic;
      spi_clk_i         : in std_logic;
      rst_i             : in std_logic;
      debug             : inout std_logic_vector(31 downto 0)
   );     
end bc_dac_ctrl;

architecture rtl of bc_dac_ctrl is

   -- wbs_bc_dac_ctrl interface:
   signal flux_fb_addr    : std_logic_vector(FLUX_FB_DAC_ADDR_WIDTH-1 downto 0);
   signal flux_fb_data    : std_logic_vector(FLUX_FB_DAC_DATA_WIDTH-1 downto 0);
   signal flux_fb_changed : std_logic;
   signal ln_bias_addr    : std_logic_vector(LN_BIAS_DAC_ADDR_WIDTH-1 downto 0);
   signal ln_bias_data    : std_logic_vector(LN_BIAS_DAC_DATA_WIDTH-1 downto 0);
   signal ln_bias_changed : std_logic;   
   
begin

   bcdc_core: bc_dac_ctrl_core
   port map(
      -- DAC hardware interface:
      flux_fb_data_o    => flux_fb_data_o,
      flux_fb_ncs_o     => flux_fb_ncs_o, 
      flux_fb_clk_o     => flux_fb_clk_o, 
      
      ln_bias_data_o    => ln_bias_data_o,
      ln_bias_ncs_o     => ln_bias_ncs_o, 
      ln_bias_clk_o     => ln_bias_clk_o, 
      
      dac_nclr_o        => dac_nclr_o,

      -- wbs_bc_dac_ctrl interface:
      flux_fb_addr_o    => flux_fb_addr,
      flux_fb_data_i    => flux_fb_data,   
      flux_fb_changed_i => flux_fb_changed,
      ln_bias_addr_o    => ln_bias_addr,
      ln_bias_data_i    => ln_bias_data,      
      ln_bias_changed_i => ln_bias_changed,   
      
      -- frame_timing signals
      update_bias_i     => update_bias_i,
      restart_frame_aligned_i => restart_frame_aligned_i,
      -- Global Signals      
      clk_i             => clk_i,
      spi_clk_i         => spi_clk_i,
      rst_i             => rst_i,
      debug             => debug
   );     
      
   -- handles wishbone transactions  
   bcdc_wbs: bc_dac_ctrl_wbs
   port map(
      -- ac_dac_ctrl interface: 32 flux_fb DACs and up to 12 low-noise bias DACs
      flux_fb_addr_i    => flux_fb_addr,
      flux_fb_data_o    => flux_fb_data,   
      flux_fb_changed_o => flux_fb_changed,
      ln_bias_addr_i    => ln_bias_addr,
      ln_bias_data_o    => ln_bias_data,      
      ln_bias_changed_o => ln_bias_changed,   
      
      -- wishbone interface:
      dat_i             => dat_i, 
      addr_i            => addr_i,
      tga_i             => tga_i, 
      we_i              => we_i,  
      stb_i             => stb_i, 
      cyc_i             => cyc_i, 
      dat_o             => dat_o, 
      ack_o             => ack_o, 

      -- global interface
      clk_i             => clk_i,
      rst_i             => rst_i,
      debug             => debug
   );
      
end rtl;