-- megafunction wizard: %ALTLVDS%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altlvds_rx 

-- ============================================================
-- File Name: adc_serdes.vhd
-- Megafunction Name(s):
-- 			altlvds_rx
--
-- Simulation Library Files(s):
-- 			altera_mf
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 8.1 Build 163 10/28/2008 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2008 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY altera_mf;
USE altera_mf.all;

ENTITY adc_serdes IS
	PORT
	(
		rx_enable		: IN STD_LOGIC  := '1';
		rx_in		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		rx_inclock		: IN STD_LOGIC  := '0';
		rx_out		: OUT STD_LOGIC_VECTOR (55 DOWNTO 0)
	);
END adc_serdes;


ARCHITECTURE SYN OF adc_serdes IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (55 DOWNTO 0);



	COMPONENT altlvds_rx
	GENERIC (
		deserialization_factor		: NATURAL;
		enable_dpa_mode		: STRING;
		implement_in_les		: STRING;
		intended_device_family		: STRING;
		lpm_hint		: STRING;
		lpm_type		: STRING;
		number_of_channels		: NATURAL;
		registered_output		: STRING;
		use_external_pll		: STRING;
		rx_align_data_reg		: STRING
	);
	PORT (
			rx_out	: OUT STD_LOGIC_VECTOR (55 DOWNTO 0);
			rx_inclock	: IN STD_LOGIC ;
			rx_in	: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
			rx_enable	: IN STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	rx_out    <= sub_wire0(55 DOWNTO 0);

	altlvds_rx_component : altlvds_rx
	GENERIC MAP (
		deserialization_factor => 7,
		enable_dpa_mode => "OFF",
		implement_in_les => "OFF",
		intended_device_family => "Stratix III",
		lpm_hint => "CBX_MODULE_PREFIX=adc_serdes",
		lpm_type => "altlvds_rx",
		number_of_channels => 8,
		registered_output => "OFF",
		use_external_pll => "ON",
		rx_align_data_reg => "RISING_EDGE"
	)
	PORT MAP (
		rx_inclock => rx_inclock,
		rx_in => rx_in,
		rx_enable => rx_enable,
		rx_out => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: Bitslip NUMERIC "7"
-- Retrieval info: PRIVATE: Channel_Data_Align_Max NUMERIC "0"
-- Retrieval info: PRIVATE: Channel_Data_Align_Reset NUMERIC "0"
-- Retrieval info: PRIVATE: Deser_Factor NUMERIC "7"
-- Retrieval info: PRIVATE: Enable_DPA_Mode STRING "OFF"
-- Retrieval info: PRIVATE: Ext_PLL STRING "ON"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix III"
-- Retrieval info: PRIVATE: Int_Device STRING "Stratix III"
-- Retrieval info: PRIVATE: LVDS_Mode NUMERIC "1"
-- Retrieval info: PRIVATE: Le_Serdes STRING "OFF"
-- Retrieval info: PRIVATE: Num_Channel NUMERIC "8"
-- Retrieval info: PRIVATE: Reg_InOut NUMERIC "0"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: Use_Data_Align NUMERIC "0"
-- Retrieval info: CONSTANT: DESERIALIZATION_FACTOR NUMERIC "7"
-- Retrieval info: CONSTANT: ENABLE_DPA_MODE STRING "OFF"
-- Retrieval info: CONSTANT: IMPLEMENT_IN_LES STRING "OFF"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix III"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "altlvds_rx"
-- Retrieval info: CONSTANT: NUMBER_OF_CHANNELS NUMERIC "8"
-- Retrieval info: CONSTANT: REGISTERED_OUTPUT STRING "OFF"
-- Retrieval info: CONSTANT: USE_EXTERNAL_PLL STRING "ON"
-- Retrieval info: CONSTANT: rx_align_data_reg STRING "RISING_EDGE"
-- Retrieval info: USED_PORT: rx_enable 0 0 0 0 INPUT VCC rx_enable
-- Retrieval info: USED_PORT: rx_in 0 0 8 0 INPUT NODEFVAL rx_in[7..0]
-- Retrieval info: USED_PORT: rx_inclock 0 0 0 0 INPUT_CLK_EXT GND rx_inclock
-- Retrieval info: USED_PORT: rx_out 0 0 56 0 OUTPUT NODEFVAL rx_out[55..0]
-- Retrieval info: CONNECT: @rx_in 0 0 8 0 rx_in 0 0 8 0
-- Retrieval info: CONNECT: rx_out 0 0 56 0 @rx_out 0 0 56 0
-- Retrieval info: CONNECT: @rx_inclock 0 0 0 0 rx_inclock 0 0 0 0
-- Retrieval info: CONNECT: @rx_enable 0 0 0 0 rx_enable 0 0 0 0
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL adc_serdes.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL adc_serdes.ppf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL adc_serdes.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL adc_serdes.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL adc_serdes.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL adc_serdes_inst.vhd FALSE
-- Retrieval info: LIB_FILE: altera_mf
-- Retrieval info: CBX_MODULE_PREFIX: ON
