-- 2003 SCUBA-2 Project
--                  All Rights Reserved

--  THIS IS UNPUBLISHED PROPRIETARY SOURCE CODE OF THE SCUBA-2 Project
--  The copyright notice above does not evidence any
--  actual or intended publication of such source code.

--  SOURCE CODE IS PROVIDED "AS IS". ALL EXPRESS OR IMPLIED CONDITIONS,
--  REPRESENTATIONS, AND WARRANTIES, INCLUDING ANY IMPLIED WARRANT OF
--  MERCHANTABILITY, SATISFACTORY QUALITY, FITNESS FOR A PARTICULAR
--  PURPOSE, OR NON-INFRINGEMENT, ARE DISCLAIMED, EXCEPT TO THE EXTENT
--  THAT SUCH DISCLAIMERS ARE HELD TO BE LEGALLY INVALID.

-- For the purposes of this code the SCUBA-2 Project consists of the
-- following organisations.

-- UKATC, Royal Observatory, Blackford Hill Edinburgh EH9 3HJ
-- UBC,   University of British Columbia, Physics & Astronomy Department,
--        Vancouver BC, V6T 1Z1

-- $Id: bc_dac_ctrl_core.vhd,v 1.13 2011-10-26 18:48:55 mandana Exp $
--
-- Project:       SCUBA2
-- Author:        Bryce Burger
-- Organisation:  UBC
--
-- Description:
-- This Blocks updates 32 + 12 serial SPI DACs on Bias Cards.
--    32 flux-fb DACs are updated simultaneously.
--    12 ln-bias DACs are updated sequentially, one after the other as
--    they share data and clock lines.
-- The flux-fb DACs are updated on every row_switch if multiplexing is on or
-- only once when new flux-fb values are written via a wishbone command
--
--
-- Revision history:
-- $Log: bc_dac_ctrl_core.vhd,v $
-- Revision 1.13  2011-10-26 18:48:55  mandana
-- chip-select is now driven by row_switch_1dly and not the spi block anymore.
-- bugfix: ln_bias is only refreshed once now, update_pending is reset at the start of the frame
-- bugfix: flux-fb is updated frame-aligned as oppose to row-aligned, this will help the internal ramp on flux-fb be synchronized on all columns.
--
-- Revision 1.12  2010/06/01 23:44:27  mandana
-- update DACs when update_bias is asserted by frame_timing instead of restart_frame
--
-- Revision 1.11  2010/05/14 22:56:10  mandana
-- all flux_fb DACs are updated at once when update_aligned is asserted
-- ln_bias lines are still updated sequentially because the data lines are shared in hardware
--
-- Revision 1.10  2010/01/28 23:29:22  mandana
-- ln_bias lines are now independently controlled.
-- the accidental bug of not driving ln_bias_data0 is now fixed!
--
-- Revision 1.9  2010/01/21 17:12:41  mandana
-- spi_clk is now generated by PLL and added to the top-level interface
-- added support for multiple ln_bias lines introduced in Bias Card Rev. E
-- parametrized flux_fb interface
-- all DACs are updated at once as oppose to sequentially
--
-- Revision 1.8  2006/04/07 22:02:21  bburger
-- Bryce:  Bug Fix:  Added integer ranges to dac_count and clk_count.  Quartus 5.1 was messing up the synthsis without these ranges.
--
-- Revision 1.7  2005/01/25 00:00:03  mandana
-- fixed the synthesis error about flux_fb_changed_reg
--
-- Revision 1.6  2005/01/20 23:08:14  mandana
-- added a register for flux_fb_changed_i
-- removed debug connections
--
-- Revision 1.5  2005/01/17 22:58:06  mandana
-- add an extra state for loading the data to the SPI module
--
-- Revision 1.4  2005/01/07 01:31:27  bench2
-- Mandana: create type dac_states
-- changed SPI modules to run at 12.5MHz
-- Now that state machine runs at 50MHz and SPI at 12.5MHz, start_spi is modified to stay high till SPI_done goes high.
-- Add an extra state NEXT_DAC2, so the dac_counter is clocked in a different state.
--
-- Revision 1.3  2005/01/04 19:19:47  bburger
-- Mandana: changed mictor assignment to 0 to 31 and swapped odd and even pods
--
-- Revision 1.2  2004/12/21 22:06:51  bburger
-- Bryce:  update
--
-- Revision 1.1  2004/11/25 03:05:08  bburger
-- Bryce:  Modified the Bias Card DAC control slaves.
--
-- Revision 1.2  2004/11/15 20:03:41  bburger
-- Bryce :  Moved frame_timing to the 'work' library, and physically moved the files to "all_cards" directory
--
-- Revision 1.1  2004/11/11 01:47:10  bburger
-- Bryce:  new
--
--   
--
-- 
-----------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
--use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library sys_param;
use sys_param.wishbone_pack.all;

library work;
use work.bias_card_pack.all;
use work.all_cards_pack.all;

entity bc_dac_ctrl_core is
   port
   (
      -- DAC hardware interface:
      -- There are 32 flux-fb DAC channels, thus 32 serial data/cs/clk lines.
      -- There are 12 (1 prior to Rev E Hardware) low-noise bias DAC channels with shared data/clk lines      
      flux_fb_data_o    : out std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);   
      flux_fb_ncs_o     : out std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);
      flux_fb_clk_o     : out std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);
      
      ln_bias_data_o    : out std_logic;                                                 -- ln_bias DAC data line (shared)
      ln_bias_ncs_o     : out std_logic_vector(NUM_LN_BIAS_DACS-1 downto 0);
      ln_bias_clk_o     : out std_logic;
      
      dac_nclr_o        : out std_logic;

      -- wbs_bc_dac_ctrl interface:
      row_addr_o        : out std_logic_vector(ROW_ADDR_WIDTH-1 downto 0);
      flux_fb_addr_o    : out std_logic_vector(FLUX_FB_DAC_ADDR_WIDTH-1 downto 0);
      flux_fb_data_i    : in flux_fb_dac_array;    
      flux_fb_changed_i : in std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);
      ln_bias_addr_o    : out std_logic_vector(LN_BIAS_DAC_ADDR_WIDTH-1 downto 0);       -- ln_bias ram address
      ln_bias_data_i    : in std_logic_vector(LN_BIAS_DAC_DATA_WIDTH-1 downto 0);        -- parallel ln_bias data
      ln_bias_changed_i : in std_logic_vector(NUM_LN_BIAS_DACS-1 downto 0);
      
      mux_flux_fb_data_i: in flux_fb_dac_array;
      enbl_mux_data_i   : in std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);
      
      -- frame_timing signals
      row_switch_i      : in std_logic;      
      update_bias_i     : in std_logic;
      restart_frame_aligned_i : in std_logic;
      restart_frame_1row_prev_i: in std_logic;
      
      -- Global Signals      
      clk_i             : in std_logic;
      spi_clk_i         : in std_logic;
      rst_i             : in std_logic;
      debug             : inout std_logic_vector(31 downto 0)
   );     
end bc_dac_ctrl_core;


architecture rtl of bc_dac_ctrl_core is
   
   -- Flux Feedback SPI interface
   signal flux_fb_data           : flux_fb_dac_array;
   signal flux_fb_dac_spi        : flux_fb_spi_array;
    
   -- Bias SPI interface
   signal ln_bias_data           : ln_bias_dac_array;
   signal ln_bias_dac_spi        : ln_bias_spi_array;
   signal ln_bias_ncs            : std_logic_vector(NUM_LN_BIAS_DACS-1 downto 0);
   signal ln_bias_ncs_1dly       : std_logic_vector(NUM_LN_BIAS_DACS-1 downto 0);
   
   -- Counter for the Flux Feedback DACs
   signal ln_bias_rd_addr        : std_logic_vector(LN_BIAS_DAC_ADDR_WIDTH-1 downto 0);             
   signal ln_bias_rd_addr_1d     : std_logic_vector(LN_BIAS_DAC_ADDR_WIDTH-1 downto 0);              -- to account for RAM read latency          
   signal row_addr               : std_logic_vector(ROW_ADDR_WIDTH-1 downto 0);
   
   -- control signals for DAC updates
   signal flux_fb_update_pending : std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);                    -- extended update-request for flux_fb
   
   signal ln_bias_dac_state      : std_logic_vector(NUM_LN_BIAS_DACS-1 downto 0);                    -- a shift register that controls which ln_bias DAC is being updated.
   signal ln_bias_update_pending : std_logic_vector(NUM_LN_BIAS_DACS-1 downto 0);                                                        -- extended frame-aligned update-request for ln_bias
   signal ln_bias_update_aligned : std_logic_vector(NUM_LN_BIAS_DACS-1 downto 0);                    -- The first ln_bias dac is updated aligned with the start of a frame and then the rest of ln_bias DACs are updated sequentially
   signal dat_rdy                : std_logic_vector(NUM_LN_BIAS_DACS-1 downto 0);
   signal ln_change_extended     : std_logic;
   
   signal update_aligned         : std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);                    -- when to update
   signal flux_fb_dat_ready      : std_logic_vector(NUM_FLUX_FB_DACS-1 downto 0);                    -- asserted all the time when multiplexing is on, otherwise, only once when flux_fb is changed
   signal row_addr_clr_pending   : std_logic;                                                        -- reset the row_address counter when a new frame has started.
   signal row_switch_1dly        : std_logic;
   
begin

   dac_nclr_o <= not rst_i;
   
   -- read-address counter for the ln-bias RAM block, note that there is 1 clock-cycle of ram latency
   ln_bias_rd_addr_counter : process (rst_i, clk_i)
   begin
      if (rst_i = '1') then
         ln_bias_rd_addr <= (others => '0');
         ln_bias_rd_addr_1d <= (others => '0');
         for i in 0 to NUM_LN_BIAS_DACS-1   loop
            ln_bias_data(i) <= x"8000"; -- mid value
         end loop;
      elsif (clk_i'event and clk_i = '1') then            
         -- if any of the values are refreshed
         if (ln_bias_update_pending(0) /= '0' or ln_bias_rd_addr = NUM_LN_BIAS_DACS-1) then  
            ln_bias_rd_addr <= (others => '0');               
         else
            ln_bias_rd_addr <= ln_bias_rd_addr + 1;       
         end if;

         ln_bias_rd_addr_1d <= ln_bias_rd_addr;
         for j in 0 to NUM_LN_BIAS_DACS-1 loop
            if (j /= conv_integer(ln_bias_rd_addr_1d)) then
               ln_bias_data(j) <= ln_bias_data(j);
            end if;   
            ln_bias_data(conv_integer(ln_bias_rd_addr_1d)) <= ln_bias_data_i;            
         end loop;
      end if;
   end process ln_bias_rd_addr_counter; 
 
   flux_fb_addr_o <= row_addr(FLUX_FB_DAC_ADDR_WIDTH-1 downto 0);
   ln_bias_addr_o <= ln_bias_rd_addr (LN_BIAS_DAC_ADDR_WIDTH-1 downto 0);

   ------------------------------------------------------------------------      
   -- delay row_switch for 1 cycle
   row_switch_1dly_proc : process (rst_i, clk_i)
   begin
      if (rst_i = '1') then
         row_switch_1dly <= '0';
      elsif (clk_i'event and clk_i = '1') then
         row_switch_1dly <= row_switch_i;
      end if;
   end process row_switch_1dly_proc;      
         
   ------------------------------------------------------------------------      
   -- row counter
   row_counter_proc : process (rst_i, clk_i)
   begin
      if (rst_i = '1') then
         row_addr <= (others =>'0');
      elsif (clk_i'event and clk_i = '1') then
         if (restart_frame_1row_prev_i = '1' and update_bias_i = '1') then 
            row_addr <= (others =>'0');
         elsif (update_bias_i = '1') then
            row_addr <= row_addr + 1;
         else
            row_addr <= row_addr;
         end if;            
      end if;
   end process row_counter_proc;      
   row_addr_o <= row_addr;
   ------------------------------------------------------------------------
   -- register previous row 
   extend_1row_prev:process(rst_i, clk_i)
   begin
     if (rst_i = '1') then
       row_addr_clr_pending <='0';
     elsif (clk_i'event and clk_i = '1') then
       if (restart_frame_1row_prev_i = '1') then
         row_addr_clr_pending <= '1';
       elsif (update_bias_i = '1') then
         row_addr_clr_pending <= '0';
       else   
         row_addr_clr_pending <= row_addr_clr_pending;
       end if;       
     end if;  
   end process; -- extend_1row_prev;
   
   ----------------------------------------------------------------------
   -- register the flux_fb change
   gen_flux_fb_update_pending: for k in 0 to NUM_FLUX_FB_DACS-1 generate
      extend_flux_fb_update:process(rst_i, clk_i)
      begin
        if (rst_i = '1') then
          flux_fb_update_pending(k) <= '0';
        elsif (clk_i'event and clk_i = '1') then
          if (flux_fb_changed_i (k) = '1') then
            flux_fb_update_pending (k) <= '1';
          elsif (update_bias_i = '1' and row_addr_clr_pending = '1') then
           flux_fb_update_pending (k) <= '0';
          else   
            flux_fb_update_pending (k) <= flux_fb_update_pending(k);
          end if;       
        end if;  
      end process; -- extend_flux_fb_update;
   end generate gen_flux_fb_update_pending;
   
   ------------------------------------------------------------------------   
   -- create ln_bias_dac_state to update the DACs
   -- since all ln_bias DACS share data and clock line, we have to update them one after the other. 
   -- hence CS of each DAC is daisy chained to next-DAC's data_rdy
   -- The first DAC, ln_bias0 is updated on the next ARZ(restart_frame_aligned)   
   ln_bias_dac_state_proc : process (rst_i, clk_i)
   begin
      if (rst_i = '1') then
         ln_bias_dac_state <= (others => '0');
         ln_bias_ncs_1dly <= (others => '0');
      elsif (clk_i'event and clk_i = '1') then
         if (restart_frame_aligned_i = '1') then 
            ln_bias_dac_state(0) <= ln_bias_update_pending(0);
         else
            ln_bias_dac_state(0) <= '0';
         end if;   
         ln_bias_ncs_1dly <= ln_bias_ncs;               
         ln_bias_dac_state(NUM_LN_BIAS_DACS-1 downto 1) <= 
                 (ln_bias_ncs_1dly(NUM_LN_BIAS_DACS-2 downto 0) xor ln_bias_ncs(NUM_LN_BIAS_DACS-2 downto 0)) and ln_bias_ncs(NUM_LN_BIAS_DACS-2 downto 0);         
      end if;
   end process ln_bias_dac_state_proc;      
   
   ------------------------------------------------------------------------   
   -- register the ln_bias change
   gen_ln_bias_update_pending: for kk in 0 to NUM_LN_BIAS_DACS-1 generate   
      extend_ln_bias_update:process(rst_i, clk_i)
      begin
      if (rst_i = '1') then
         ln_bias_update_pending(kk) <= '0';       
      elsif (clk_i'event and clk_i = '1') then
        if (ln_bias_dac_state(kk) = '1') then
            ln_bias_update_pending(kk) <= '0';
         elsif (ln_bias_changed_i(kk) = '1') then
            ln_bias_update_pending(kk) <= '1';
         else   
            ln_bias_update_pending(kk) <= ln_bias_update_pending(kk);
         end if;       
      end if;  
      end process; -- extend_ln_bias_update_all;
   end generate;   
      
   ln_bias_update_aligned(NUM_LN_BIAS_DACS-1 downto 0) <= (others => '1');
   
   ------------------------------------------------------------------------
   -- Instantiate spi interface blocks for flux-fb dacs
   gen_spi_flux_fb: for k in 0 to NUM_FLUX_FB_DACS-1 generate
      -- flux-fb DACs are refreshed:
      -- on every row_switch when multiplexing is on (enbl_mux = 1)
      -- only when new values are written (through wishbone interface) when multiplexing is off (enbl_mux = 0) 
      update_aligned(k) <= update_bias_i when enbl_mux_data_i(k) = '1' else
                           (restart_frame_aligned_i and flux_fb_update_pending(k));
      
      flux_fb_dat_ready(k) <= enbl_mux_data_i(k) or flux_fb_changed_i(k); 
      
      flux_fb_data(k) <= mux_flux_fb_data_i(k) when enbl_mux_data_i(k) = '1' else 
                              flux_fb_data_i(k);
                      
      spi_dac_ctrl_i: spi_dac_ctrl
      generic map (
         DAC_DATA_WIDTH      => FLUX_FB_DAC_DATA_WIDTH
      )   
      port map (  
         -- global signals
         rst_i               => rst_i,
         clk_25_i            => spi_clk_i,
         clk_50_i            => clk_i,
              
         -- control signals from frame timing block
         restart_frame_aligned_i => update_aligned(k),
         
         -- control signal indicates dat_i is updated
         dat_rdy_i           => flux_fb_dat_ready(k) ,
         
         -- parallel data to be serialized
         dat_i               => flux_fb_data(k), 
         
         -- SPI interface to MAX 5443 DAC
         dac_spi_o           => flux_fb_dac_spi (k)
      );   
      -- Bit 2:  chip select (active low)
      -- Bit 1:  serial clock out
      -- Bit 0:  serial data out
      flux_fb_ncs_o (k)  <= flux_fb_dac_spi(k)(2) when enbl_mux_data_i(k) = '0' else row_switch_1dly;
      flux_fb_clk_o (k)  <= flux_fb_dac_spi(k)(1);
      flux_fb_data_o (k) <= flux_fb_dac_spi(k)(0) when rst_i ='0' else '0';
      
   end generate gen_spi_flux_fb;
   
   ------------------------------------------------------------------------
   -- Instantiate spi interface blocks for ln_bias dacs
   ------------------------------------------------------------------------
   gen_spi_ln_bias: for k in 0 to NUM_LN_BIAS_DACS-1 generate
      
      dat_rdy(k) <= ln_bias_dac_state(k) and ln_bias_update_pending(k);
      
      spi_dac_ctrl_i: spi_dac_ctrl
      generic map (
         DAC_DATA_WIDTH      => LN_BIAS_DAC_DATA_WIDTH
      )   
      port map (  
         -- global signals
         rst_i               => rst_i,
         clk_25_i            => spi_clk_i,
         clk_50_i            => clk_i,
              
         -- control signals from frame timing block
         restart_frame_aligned_i => ln_bias_update_aligned(k),
         
         -- control signal indicates dat_i is updated
         dat_rdy_i           => dat_rdy(k), 
         
         -- parallel data to be serialized
         dat_i               => ln_bias_data(k), 
         
         -- SPI interface to MAX 5443 DAC
         dac_spi_o           => ln_bias_dac_spi (k)
      );   
      -- Bit 2:  chip select (active low)
      -- Bit 1:  serial clock out
      -- Bit 0:  serial data out
      ln_bias_ncs_o (k)  <= ln_bias_dac_spi(k)(2) when rst_i = '0' else '1';
      ln_bias_ncs (k) <= ln_bias_dac_spi(k)(2); 
--      ln_bias_clk_o (k)  <= ln_bias_dac_spi(k)(1);
--      ln_bias_data_o (k) <= ln_bias_dac_spi(k)(0);
            
   end generate gen_spi_ln_bias;
   ln_bias_clk_o  <= ln_bias_dac_spi(11)(1) or ln_bias_dac_spi(10)(1) or ln_bias_dac_spi(9)(1) or ln_bias_dac_spi(8)(1) or
                     ln_bias_dac_spi(7)(1) or ln_bias_dac_spi(6)(1) or ln_bias_dac_spi(5)(1) or ln_bias_dac_spi(4)(1) or
                     ln_bias_dac_spi(3)(1) or ln_bias_dac_spi(2)(1) or ln_bias_dac_spi(1)(1) or ln_bias_dac_spi(0)(1);
   ln_bias_data_o <= ln_bias_dac_spi(11)(0) or ln_bias_dac_spi(10)(0) or ln_bias_dac_spi(9)(0) or ln_bias_dac_spi(8)(0) or
                     ln_bias_dac_spi(7)(0) or ln_bias_dac_spi(6)(0) or ln_bias_dac_spi(5)(0) or ln_bias_dac_spi(4)(0) or
                     ln_bias_dac_spi(3)(0) or ln_bias_dac_spi(2)(0) or ln_bias_dac_spi(1)(0) or ln_bias_dac_spi(0)(0); 
                     
end rtl;