-- Copyright (c) 2003 SCUBA-2 Project
--               All Rights Reserved
--
-- THIS IS UNPUBLISHED PROPRIETARY SOURCE CODE OF THE SCUBA-2 Project
-- The copyright notice above does not evidence any
-- actual or intended publication of such source code.
--
-- SOURCE CODE IS PROVIDED "AS IS". ALL EXPRESS OR IMPLIED CONDITIONS,
-- REPRESENTATIONS, AND WARRANTIES, INCLUDING ANY IMPLIED WARRANT OF
-- MERCHANTABILITY, SATISFACTORY QUALITY, FITNESS FOR A PARTICULAR
-- PURPOSE, OR NON-INFRINGEMENT, ARE DISCLAIMED, EXCEPT TO THE EXTENT
-- THAT SUCH DISCLAIMERS ARE HELD TO BE LEGALLY INVALID.
--
-- For the purposes of this code the SCUBA-2 Project consists of the
-- following organisations.
--
-- UKATC, Royal Observatory, Blackford Hill Edinburgh EH9 3HJ
-- UBC,   University of British Columbia, Physics & Astronomy Department,
--        Vancouver BC, V6T 1Z1
--
-- $Id: cmd_queue.vhd,v 1.20 2004/07/16 18:23:20 erniel Exp $
--
-- Project:    SCUBA2
-- Author:     Bryce Burger
-- Organisation:  UBC
--
-- Description:
-- This file implements the cmd_queue block in the issue/reply hardware
-- on the clock card.
--
-- Revision history:
-- $Log: cmd_queue.vhd,v $
-- Revision 1.20  2004/07/16 18:23:20  erniel
-- in progress
--
-- Revision 1.19  2004/07/07 00:35:23  bburger
-- in progress
--
-- Revision 1.18  2004/06/30 23:10:53  bburger
-- in progress
--
-- Revision 1.17  2004/06/19 01:16:13  bburger
-- send fsm bug fixes
--
-- Revision 1.16  2004/06/16 17:02:36  bburger
-- in progress
--
-- Revision 1.1  2004/05/11 02:17:31  bburger
-- new
--
--
------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library sys_param;
use sys_param.wishbone_pack.all;
use sys_param.frame_timing_pack.all;

library components;
use components.component_pack.all;

library work;
use work.issue_reply_pack.all;
use work.cmd_queue_ram40_pack.all;
use work.async_pack.all;

entity cmd_queue is
   port(
      -- reply_queue interface
      uop_status_i  : in std_logic_vector(UOP_STATUS_BUS_WIDTH-1 downto 0); -- Tells the cmd_queue whether a reply was successful or erroneous
      uop_rdy_o     : out std_logic; -- Tells the reply_queue when valid m-op and u-op codes are asserted on it's interface
      uop_ack_i     : in std_logic; -- Tells the cmd_queue that a reply to the u-op waiting to be retired has been found and it's status is asserted on uop_status_i
      uop_discard_o : out std_logic; -- Tells the reply_queue whether or not to discard the reply to the current u-op reply when uop_rdy_i goes low.  uop_rdy_o can only go low after rq_ack_o has been received.
      uop_timedout_o: out std_logic; -- Tells that reply_queue that it should generated a timed-out reply based on the the par_id, card_addr, etc of the u-op being retired.
      uop_o         : out std_logic_vector(QUEUE_WIDTH-1 downto 0); --Tells the reply_queue the next u-op that the cmd_queue wants to retire

      -- cmd_translator interface
      card_addr_i   : in std_logic_vector (CARD_ADDR_BUS_WIDTH-1 downto 0); -- The card address of the m-op
      par_id_i      : in std_logic_vector (PAR_ID_BUS_WIDTH-1 downto 0); -- The parameter id of the m-op
      data_size_i   : in std_logic_vector (DATA_SIZE_BUS_WIDTH-1 downto 0); -- The number of 32-bit words of data in the m-op
      data_i        : in std_logic_vector (DATA_BUS_WIDTH-1 downto 0);  -- Data belonging to a m-op
      data_clk_i    : in std_logic; -- Clocks in 32-bit wide data
      mop_i         : in std_logic_vector (MOP_BUS_WIDTH-1 downto 0); -- M-op sequence number
      issue_sync_i  : in std_logic_vector (SYNC_NUM_BUS_WIDTH-1 downto 0); -- The issuing sync-pulse sequence number
      mop_rdy_i     : in std_logic; -- Tells cmd_queue when a m-op is ready
      mop_ack_o     : out std_logic; -- Tells the cmd_translator when cmd_queue has taken the m-op and is ready to receive data
      
      -- lvds_tx interface
      tx_o          : out std_logic;  -- transmitter output pin
      clk_25mhz_i   : in std_logic;  -- PLL locked 25MHz input clock for the

      -- Clock lines
      sync_i        : in std_logic; -- The sync pulse determines when and when not to issue u-ops
      clk_i         : in std_logic; -- Advances the state machines
      clk_400mhz_i  : in std_logic; -- Fast clock used for doing multi-cycle operations (inserting and deleting u-ops from the command queue) in a single clk_i cycle.  clk_400mhz_i must be at least 2x as fast as clk_i
      rst_i         : in std_logic  -- Resets all FSMs
   );
end cmd_queue;

architecture behav of cmd_queue is

constant ADDR_ZERO          : std_logic_vector(QUEUE_ADDR_WIDTH-1 downto 0) := (others => '0');
constant ADDR_FULL_SCALE    : std_logic_vector(QUEUE_ADDR_WIDTH-1 downto 0) := (others => '1');
constant TIMEOUT_LEN        : std_logic_vector(TIMEOUT_SYNC_BUS_WIDTH-1 downto 0) := "00000001";  -- The number of sync pulses after which an instruction will expire
constant MAX_SYNC_COUNT     : integer := 255;

-- Command queue inputs/ouputs (this interface was generated by a Quartus II megafunction for a RAM block)
signal data_sig             : std_logic_vector(QUEUE_WIDTH-1 downto 0);
signal wraddress_sig        : std_logic_vector(7 downto 0);
signal rdaddress_a_sig      : std_logic_vector(7 downto 0);
signal rdaddress_b_sig      : std_logic_vector(7 downto 0);
signal wren_sig             : std_logic;
signal qa_sig               : std_logic_vector(QUEUE_WIDTH-1 downto 0);
signal qb_sig               : std_logic_vector(QUEUE_WIDTH-1 downto 0);
signal nfast_clk            : std_logic;
signal n_clk                : std_logic;

-- Indicates the number u-ops contained in the command queue
signal uop_counter          : std_logic_vector(UOP_BUS_WIDTH - 1 downto 0);

-- Sync-pulse counter inputs/outputs.  These are used to determine when u-ops have expired.
signal sync_count_slv       : std_logic_vector(7 downto 0);
signal sync_count_int       : integer;
signal clk_count            : integer;
signal clk_error            : std_logic_vector(31 downto 0);

-- Command queue management variables
signal uops_generated       : integer;
signal cards_addressed      : integer;
signal num_uops             : integer;
signal data_size_int        : integer;
signal size_uops            : integer;
-- num_uops_inserted:  determines when to stop inserting u-ops
signal num_uops_inserted    : integer;
signal queue_space          : integer := QUEUE_LEN;

-- Command queue address pointers.  Each one of these are managed by a different FSM.
signal retire_ptr           : std_logic_vector(QUEUE_ADDR_WIDTH-1 downto 0);
signal flush_ptr            : std_logic_vector(QUEUE_ADDR_WIDTH-1 downto 0);
signal send_ptr             : std_logic_vector(QUEUE_ADDR_WIDTH-1 downto 0);
signal free_ptr             : std_logic_vector(QUEUE_ADDR_WIDTH-1 downto 0);

-- Insertion FSM:  inserts u-ops into the command queue
type insert_states is (IDLE, INSERT_HDR1, INSERT_HDR2, INSERT_DATA, DONE, RESET, STALL);
signal present_insert_state : insert_states;
signal next_insert_state    : insert_states;
signal data_count           : std_logic_vector(CQ_DATA_SIZE_BUS_WIDTH-1 downto 0);
-- insert_uop_ack:  tells the generate FSM when the insert FSM is ready to insert the next u-op
signal insert_uop_ack       : std_logic;
-- inserting:  used to keep track of how much space there is in the queue.
-- To keep track of space, it is asserted until the insert FSM asserts finishes inserting a u-op
signal inserting            : std_logic;

-- Retire FSM:  waits for replies from the Bus Backplane, and retires pending instructions in the the command queue
type retire_states is (IDLE, NEXT_UOP, STATUS, RETIRE, FLUSH, EJECT, NEXT_FLUSH, FLUSH_STATUS, RESET);
signal present_retire_state : retire_states;
signal next_retire_state    : retire_states;
signal retired              : std_logic; --Out, to the u-op counter fsm
signal uop_timed_out        : std_logic;

-- Generate FSM:  translates M-ops into u-ops
type gen_uop_states is (IDLE, INSERT, PS_CARD, CLOCK_CARD, ADDR_CARD, READOUT_CARD1, READOUT_CARD2, READOUT_CARD3, READOUT_CARD4, BIAS_CARD1, BIAS_CARD2, BIAS_CARD3, CLEANUP, RESET, DONE);
signal present_gen_state    : gen_uop_states;
signal next_gen_state       : gen_uop_states;
signal new_insert_state     : gen_uop_states;
signal mop_rdy              : std_logic; --In from the previous block in the chain
-- insert_uop_rdy:  tells the insert FSM when a new u-op is available
signal insert_uop_rdy       : std_logic; --Out, to insertion fsm
signal new_card_addr        : std_logic_vector(CQ_CARD_ADDR_BUS_WIDTH-1 downto 0); --out, to insertion fsm
signal new_par_id           : std_logic_vector(CQ_PAR_ID_BUS_WIDTH-1 downto 0) := x"00"; --out, to insertion fsm.  This is a hack.

-- Send FSM:  sends u-ops over the bus backplane
type send_states is (LOAD, ISSUE, HEADER_A, HEADER_B, DATA, CHECKSUM, NEXT_UOP, RESET);
signal present_send_state   : send_states;
signal next_send_state      : send_states;
-- This signal needs support in the send FSM.  So far I have not implemented this.
signal freeze_send          : std_logic;  --In, freezes the send pointer when flushing out invalidated u-ops
signal uop_send_expired     : std_logic;
signal issue_sync           : std_logic_vector (SYNC_NUM_BUS_WIDTH-1 downto 0);
signal timeout_sync         : std_logic_vector (SYNC_NUM_BUS_WIDTH-1 downto 0);

-- Wishbone signals to/from async_tx
signal cmd_tx_dat           : std_logic_vector (31 downto 0);
signal cmd_tx_start         : std_logic;
signal cmd_tx_done          : std_logic;

-- CRC signals:
signal crc_clr              : std_logic;
signal crc_num_bits         : integer;
signal crc_data             : std_logic;
signal crc_done             : std_logic;
signal crc_valid            : std_logic;
signal crc_checksum         : std_logic_vector(CHECKSUM_BUS_WIDTH-1 downto 0);

-- Constants that can be removed when the sync_counter and frame_timer are moved out of this block
constant HIGH               : std_logic := '1';
constant LOW                : std_logic := '0';
constant INT_ZERO           : integer := 0;

begin
   -- Command queue (FIFO)
   cmd_queue_ram40_inst: cmd_queue_ram40_test
      port map(
         data        => data_sig,
         wraddress   => wraddress_sig,
         rdaddress_a => rdaddress_a_sig,
         rdaddress_b => rdaddress_b_sig,
         wren        => wren_sig,
         clock       => n_clk,
         -- qa_sig data are used by the send FSM
         qa          => qa_sig,
         -- qb_sig data are used by the retire FSM
         qb          => qb_sig
      );

   -- The sync counter will be moved outside this block
   sync_counter: counter
      generic map(MAX => MAX_SYNC_COUNT)
      port map(
         clk_i       => sync_i,
         rst_i       => rst_i,
         ena_i       => HIGH,
         load_i      => LOW,
         down_i      => LOW,
         count_i     => INT_ZERO,
         count_o     => sync_count_int
      );

   frame_timer: frame_timing
     port map(
         clk_i       => clk_i,
         sync_i      => sync_i,
         frame_rst_i => rst_i,
         clk_count_o => clk_count,
         clk_error_o => clk_error
     );

   -- lvds_tx is the LVDS interface to the Bus Backplane
   cmd_tx: lvds_tx
      port map(
         clk_i      => clk_i,
         comm_clk_i => clk_25mhz_i,
         rst_i      => rst_i,
         dat_i      => cmd_tx_dat,
         start_i    => cmd_tx_start,
         done_o     => cmd_tx_done,
         lvds_o     => tx_o
      );
      
   cmd_crc: crc
      generic map(
         POLY_WIDTH  => CHECKSUM_BUS_WIDTH
      )
      port map(
         clk        => clk_25mhz_i,
         rst        => rst_i,
         clr_i      => crc_clr,
         ena_i      => '1',
         data_i     => crc_data,
         num_bits_i => crc_num_bits,
         poly_i     => "00000100110000010001110110110111",  --CRC-32        
         done_o     => crc_done,
         valid_o    => crc_valid,
         checksum_o => crc_checksum 
      );

   -- Counter for tracking free space in the queue:
   space_calc: process(clk_i, rst_i)
   begin
      if(rst_i = '1') then
         queue_space <= QUEUE_LEN;
      elsif(clk_i'event and clk_i = '1') then
         if(inserting = '1' and retired = '0') then
            queue_space <= queue_space - 1;
         elsif(inserting = '0' and retired = '1') then
            queue_space <= queue_space + 1;
         -- All other operations balance each other out
         end if;
      end if;
   end process;

   -- FSM for inserting u-ops into the u-op queue
   -- Assumes that clk_400mhz_i is in phase with clk_i
   insert_state_FF: process(clk_i, rst_i)
   begin
      if(rst_i = '1') then
         present_insert_state <= RESET;
      elsif(clk_i'event and clk_i = '1') then
         present_insert_state <= next_insert_state;
      end if;
   end process;

   insert_state_NS: process(present_insert_state, insert_uop_rdy, present_gen_state)
   begin
      case present_insert_state is
         when RESET =>
            next_insert_state <= IDLE;
         when IDLE =>
            -- The gen_state FSM will only try to add a u-op to the queue if there is space available, so no checking is necessary here.
            -- ***This needs to react as soon as there is a u-op ready to insert..
            if(insert_uop_rdy = '1') then
               next_insert_state <= INSERT_HDR1;
            else
               next_insert_state <= IDLE;
            end if;
         when INSERT_HDR1 =>
            next_insert_state <= INSERT_HDR2;
         when INSERT_HDR2 =>
            if(data_size_i(CQ_DATA_SIZE_BUS_WIDTH-1 downto 0) = x"0000") then
               next_insert_state <= DONE;
            else
               next_insert_state <= INSERT_DATA;
            end if;
         when INSERT_DATA =>
            -- INSERT_DATA state has to loop without any others in between to make sure that it records all data from the cmd_translator block
            if(data_count < data_size_i(CQ_DATA_SIZE_BUS_WIDTH-1 downto 0)) then
               next_insert_state <= INSERT_DATA;
            else
               next_insert_state <= DONE;
            end if;
         when DONE =>
            next_insert_state <= STALL;
         -- This state exists to delay the FSM from returning too quickly to the IDLE state and trying to insert the same u-op again.
         -- The side effect of this state is that the u-op is only inserted on the second clk_400mhz_i cycle after it becomes available for insertion
         when STALL =>
            if(new_insert_state /= present_gen_state and
              (present_gen_state = PS_CARD or
               present_gen_state = CLOCK_CARD or
               present_gen_state = ADDR_CARD or
               present_gen_state = READOUT_CARD1 or
               present_gen_state = READOUT_CARD2 or
               present_gen_state = READOUT_CARD3 or
               present_gen_state = READOUT_CARD4 or
               present_gen_state = BIAS_CARD1 or
               present_gen_state = BIAS_CARD2 or
               present_gen_state = BIAS_CARD3)) then
               next_insert_state <= IDLE;
            else
               next_insert_state <= STALL;
            end if;
         when others =>
            next_insert_state <= IDLE;
      end case;
   end process;

   insert_state_out: process(present_insert_state, mop_i, uop_counter, issue_sync_i, new_card_addr, new_par_id, present_gen_state)
   -- There is something sketchy about the sensitivity list.  free_ptr does not appear anywhere on the list.  It can't because of my free_ptr <= free_ptr + 1 statement below.  However, it should because it appears on the lhs in the INSERT state
   begin
      case present_insert_state is
         when RESET =>
            wren_sig       <= '0';
            data_count     <= x"0000";
            mop_ack_o      <= '0';
            insert_uop_ack <= '0';
            free_ptr       <= ADDR_ZERO;
            inserting      <= '0';
         when IDLE =>
            -- The RAM block and the functions that write to it will be operating at higher speed than the rest of the logic.
            -- INSERT and DONE should complete in less than one clk_i cycle for this to work
            wren_sig       <= '0';
            data_count     <= x"0000";
            mop_ack_o      <= '0';
            insert_uop_ack <= '0';
            inserting      <= '0';
         when INSERT_HDR1 =>
            wren_sig       <= '1';
            data_count     <= x"0000";
            mop_ack_o      <= '0';
            insert_uop_ack <= '0';
            inserting      <= '1';
            data_sig(QUEUE_WIDTH-1      downto ISSUE_SYNC_END)   <= issue_sync_i;
            data_sig(ISSUE_SYNC_END-1   downto TIMEOUT_SYNC_END) <= issue_sync_i + TIMEOUT_LEN;
            data_sig(TIMEOUT_SYNC_END-1 downto DATA_SIZE_END)    <= data_size_i(CQ_DATA_SIZE_BUS_WIDTH-1 downto 0);
            wraddress_sig <= free_ptr;
         when INSERT_HDR2 =>
            wren_sig       <= '1';
            data_count     <= x"0000";
            mop_ack_o      <= '1';
            insert_uop_ack <= '0';
            inserting      <= '1';
            -- In this state, I need to assert the 
            data_sig(QUEUE_WIDTH-1      downto CARD_ADDR_END)    <= new_card_addr;
            data_sig(CARD_ADDR_END-1    downto PARAM_ID_END)     <= new_par_id;
            data_sig(PARAM_ID_END-1     downto MOP_END)          <= mop_i;
            -- new u-op sequence number.  This FSM automatically increments uop_counter after a u-op is added.
            data_sig(MOP_END-1          downto UOP_END)          <= uop_counter;
            wraddress_sig <= free_ptr;
            -- After adding new u-op header1 info:
            if(free_ptr = ADDR_FULL_SCALE) then
               free_ptr <= ADDR_ZERO;
            else
               free_ptr <= free_ptr + 1;
            end if;
         when INSERT_DATA =>
            wren_sig       <= '1';
            data_count     <= data_count + 1;
            mop_ack_o      <= '0';
            insert_uop_ack <= '0';
            inserting      <= '1';
            wraddress_sig <= free_ptr;
            if(next_insert_state = DONE) then
               -- This is here so that the STALL state can detect when the Generate FSM tries to issue a new u-op
               -- The Insert FSM will remain stalled until it detetects a new u-op from the Generate FSM
               new_insert_state <= present_gen_state;
            end if;
            -- After adding new u-op header2 info, or data:
            if(free_ptr = ADDR_FULL_SCALE) then
               free_ptr <= ADDR_ZERO;
            else
               free_ptr <= free_ptr + 1;
            end if;
         when DONE =>
            wren_sig       <= '0';
            data_count     <= x"0000";
            mop_ack_o      <= '0';
            insert_uop_ack <= '1';
            inserting      <= '0';
            -- After adding a new u-op:
            if(free_ptr = ADDR_FULL_SCALE) then
               free_ptr <= ADDR_ZERO;
            else
               free_ptr <= free_ptr + 1;
            end if;
         when STALL =>
            wren_sig       <= '0';
            data_count     <= x"0000";
            mop_ack_o      <= '0';
            insert_uop_ack <= '0';
            inserting      <= '0';
         when others =>
            wren_sig       <= '0';
            data_count     <= x"0000";
            mop_ack_o      <= '0';
            insert_uop_ack <= '0';
            inserting      <= '0';
      end case;
   end process;

   -- Retire FSM:
   retire_state_FF: process(clk_i, rst_i)
   begin
      if(rst_i = '1') then
         present_retire_state <= RESET;
      elsif(clk_i'event and clk_i = '1') then
         present_retire_state <= next_retire_state;
      end if;
   end process retire_state_FF;

   uop_timed_out <= '1' when (sync_count_slv > qb_sig(ISSUE_SYNC_END - 1 downto TIMEOUT_SYNC_END) or
                             (sync_count_slv < qb_sig(ISSUE_SYNC_END - 1 downto TIMEOUT_SYNC_END) and MAX_SYNC_COUNT - qb_sig(ISSUE_SYNC_END - 1 downto TIMEOUT_SYNC_END) + sync_count_slv > TIMEOUT_LEN)) else '0';

   retire_state_NS: process(present_retire_state, retire_ptr, send_ptr, uop_ack_i, uop_status_i, uop_timed_out)
   begin
      case present_retire_state is
         when RESET =>
            next_retire_state <= IDLE;
         when IDLE =>
            if(retire_ptr /= send_ptr) then
               next_retire_state <= NEXT_UOP;
            else
               next_retire_state <= IDLE;
            end if;
         when NEXT_UOP =>
            next_retire_state <= STATUS;
         when STATUS =>
            if(uop_ack_i = '1') then
               if(uop_status_i = SUCCESS) then
                  next_retire_state <= RETIRE;
               elsif(uop_status_i = FAIL) then
                  next_retire_state <= FLUSH;
               --Instruction timed out
               elsif(uop_timed_out = '1') then
                  next_retire_state <= EJECT;
               end if;
            elsif (uop_ack_i = '0') then
               next_retire_state <= STATUS;
            end if;
         when RETIRE =>
            next_retire_state <= IDLE;
         when FLUSH =>
            if(retire_ptr /= send_ptr) then
               next_retire_state <= NEXT_FLUSH;
            elsif(retire_ptr = send_ptr) then
               next_retire_state <= IDLE;
            end if;
         when EJECT =>
            next_retire_state <= IDLE;
         when NEXT_FLUSH =>
            next_retire_state <= FLUSH_STATUS;
         when FLUSH_STATUS =>
            if(uop_ack_i = '0') then
               next_retire_state <= FLUSH_STATUS;
            elsif(uop_ack_i = '1') then
               next_retire_state <= FLUSH;
            end if;
         when others =>
            next_retire_state <= IDLE;
      end case;
   end process;

   rdaddress_b_sig <= retire_ptr;
   uop_o <= qb_sig;

   retire_state_out: process(present_retire_state)
   begin
      case present_retire_state is
         when RESET =>
            uop_rdy_o      <= '0';
            freeze_send    <= '0';
            uop_timedout_o <= '0';
            uop_discard_o  <= '0';
            retire_ptr     <= ADDR_ZERO;
            flush_ptr      <= ADDR_ZERO;
            retired        <= '0';
         when IDLE =>
            uop_rdy_o      <= '0';
            freeze_send    <= '0';
            uop_timedout_o <= '0';
            uop_discard_o  <= '0';
            retired        <= '0';
         when NEXT_UOP =>
            uop_rdy_o      <= '1';
            freeze_send    <= '0';
            uop_timedout_o <= '0';
            uop_discard_o  <= '0';
            retired        <= '0';
         when STATUS =>
            uop_rdy_o      <= '1';
            freeze_send    <= '0';
            uop_timedout_o <= '0';
            uop_discard_o  <= '0';
            retired        <= '0';
         when RETIRE =>
            uop_rdy_o      <= '0';
            freeze_send    <= '0';
            uop_timedout_o <= '0';
            uop_discard_o  <= '0';
            retired        <= '1';
            retire_ptr     <= retire_ptr + 2 + qb_sig(DATA_SIZE_END+QUEUE_ADDR_WIDTH-1 downto DATA_SIZE_END);
            flush_ptr      <= flush_ptr + 2 + qb_sig(DATA_SIZE_END+QUEUE_ADDR_WIDTH-1 downto DATA_SIZE_END);
         when FLUSH =>
            uop_rdy_o      <= '0';
            freeze_send    <= '1';
            uop_timedout_o <= '0';
            uop_discard_o  <= '1';
            retired        <= '1';
         when EJECT =>
            uop_rdy_o      <= '0';
            freeze_send    <= '0';
            uop_timedout_o <= '1';
            uop_discard_o  <= '1';
            retired        <= '1';
            retire_ptr     <= retire_ptr + 2 + qb_sig(DATA_SIZE_END+QUEUE_ADDR_WIDTH-1 downto DATA_SIZE_END);
            flush_ptr      <= flush_ptr + 2 + qb_sig(DATA_SIZE_END+QUEUE_ADDR_WIDTH-1 downto DATA_SIZE_END);
         when NEXT_FLUSH =>
            uop_rdy_o      <= '1';
            freeze_send    <= '1';
            uop_timedout_o <= '0';
            uop_discard_o  <= '1';
            retired        <= '0';
            flush_ptr      <= flush_ptr + 2 + qb_sig(DATA_SIZE_END+QUEUE_ADDR_WIDTH-1 downto DATA_SIZE_END);
         when FLUSH_STATUS =>
            uop_rdy_o      <= '1';
            freeze_send    <= '1';
            uop_timedout_o <= '0';
            uop_discard_o  <= '1';
            retired        <= '0';
         when others =>
            uop_rdy_o      <= '0';
            freeze_send    <= '0';
            uop_timedout_o <= '0';
            uop_discard_o  <= '0';
            retired        <= '0';
      end case;
   end process;

   -- Generate FSM:
   gen_state_FF: process(clk_i, rst_i)
   begin
      if(rst_i = '1') then
         present_gen_state <= RESET;
      elsif(clk_i'event and clk_i = '1') then
         present_gen_state <= next_gen_state;
      end if;
   end process;

   gen_state_NS: process(present_gen_state, mop_rdy, queue_space, num_uops, par_id_i, card_addr_i, new_par_id, size_uops)
   begin
      case present_gen_state is
         when RESET =>
            next_gen_state <= IDLE;
         when IDLE =>
            if(mop_rdy = '0') then
               next_gen_state <= IDLE;
            elsif(mop_rdy = '1') then
               if(queue_space < size_uops) then
                  next_gen_state <= IDLE;
               elsif(queue_space >= size_uops) then
                  next_gen_state <= INSERT;
               end if;
            end if;
         when INSERT =>
            if(card_addr_i = BCS) then
               next_gen_state <= BIAS_CARD1;
            elsif(card_addr_i = RCS) then
               next_gen_state <= READOUT_CARD1;
            elsif(card_addr_i = ALL_FBGA_CARDS) then
               next_gen_state <= ADDR_CARD;
            elsif(card_addr_i = ALL_CARDS) then
               next_gen_state <= PS_CARD;
            elsif(card_addr_i = PSC) then
               next_gen_state <= PS_CARD;
            elsif(card_addr_i = CC) then
               next_gen_state <= CLOCK_CARD;
            elsif(card_addr_i = AC) then
               next_gen_state <= ADDR_CARD;
            elsif(card_addr_i = RC1) then
               next_gen_state <= READOUT_CARD1;
            elsif(card_addr_i = RC2) then
               next_gen_state <= READOUT_CARD2;
            elsif(card_addr_i = RC3) then
               next_gen_state <= READOUT_CARD3;
            elsif(card_addr_i = RC4) then
               next_gen_state <= READOUT_CARD4;
            elsif(card_addr_i = BC1) then
               next_gen_state <= BIAS_CARD1;
            elsif(card_addr_i = BC2) then
               next_gen_state <= BIAS_CARD2;
            elsif(card_addr_i = BC3) then
               next_gen_state <= BIAS_CARD3;
            else
               next_gen_state <= CLEANUP;  -- Catch all invalid card_id's with this statement
            end if;
         when PS_CARD =>
            if(card_addr_i = ALL_CARDS) then
               next_gen_state <= CLOCK_CARD;
            elsif(card_addr_i = PSC) then
               next_gen_state <= CLEANUP;
            end if;
         when CLOCK_CARD =>
            if(card_addr_i = ALL_CARDS or card_addr_i = ALL_FBGA_CARDS) then
               next_gen_state <= ADDR_CARD;
            elsif(card_addr_i = CC) then
               next_gen_state <= CLEANUP;
            end if;
         when ADDR_CARD =>
            if(card_addr_i = ALL_CARDS or card_addr_i = ALL_FBGA_CARDS) then
               next_gen_state <= READOUT_CARD1;
            elsif(card_addr_i = AC) then
               next_gen_state <= CLEANUP;
            end if;
         when READOUT_CARD1 =>
            if(card_addr_i = ALL_CARDS or card_addr_i = ALL_FBGA_CARDS or card_addr_i = RCS) then
               next_gen_state <= READOUT_CARD2;
            elsif(card_addr_i = RC1) then
               next_gen_state <= CLEANUP;
            end if;
         when READOUT_CARD2 =>
            if(card_addr_i = ALL_CARDS or card_addr_i = ALL_FBGA_CARDS or card_addr_i = RCS) then
               next_gen_state <= READOUT_CARD3;
            elsif(card_addr_i = RC2) then
               next_gen_state <= CLEANUP;
            end if;
         when READOUT_CARD3 =>
            if(card_addr_i = ALL_CARDS or card_addr_i = ALL_FBGA_CARDS or card_addr_i = RCS) then
               next_gen_state <= READOUT_CARD4;
            elsif(card_addr_i = RC3) then
               next_gen_state <= CLEANUP;
            end if;
         when READOUT_CARD4 =>
            if(card_addr_i = ALL_CARDS or card_addr_i = ALL_FBGA_CARDS) then
               next_gen_state <= BIAS_CARD1;
            elsif(card_addr_i = RC4 or card_addr_i = RCS) then
               next_gen_state <= CLEANUP;
            end if;
         when BIAS_CARD1 =>
            if(card_addr_i = ALL_CARDS or card_addr_i = ALL_FBGA_CARDS or card_addr_i = BCS) then
               next_gen_state <= BIAS_CARD2;
            elsif(card_addr_i = BC1) then
               next_gen_state <= CLEANUP;
            end if;
         when BIAS_CARD2 =>
            if(card_addr_i = ALL_CARDS or card_addr_i = ALL_FBGA_CARDS or card_addr_i = BCS) then
               next_gen_state <= BIAS_CARD3;
            elsif(card_addr_i = BC2) then
               next_gen_state <= CLEANUP;
            end if;
         when BIAS_CARD3 =>
            if(card_addr_i = ALL_CARDS or card_addr_i = ALL_FBGA_CARDS) then
               next_gen_state <= CLEANUP;
            elsif(card_addr_i = BC3 or card_addr_i = BCS) then
               next_gen_state <= CLEANUP;
            end if;
         when CLEANUP =>
            if(insert_uop_ack = '1') then
               -- Monitor all the exit points from this sequence of states.
               if(par_id_i(7 downto 0) = RET_DAT_ADDR or par_id_i(7 downto 0) = STATUS_ADDR) then
                  -- CYC_OO_SYNC is the last u-op instruction in a RET_DAT or STATUS m-op.
                  -- RET_DAT and STATUS are the only m-op that generate u-ops with different command codes
                  if(num_uops_inserted /= num_uops) then
                     if(card_addr_i = BCS) then
                        next_gen_state <= BIAS_CARD1;
                     elsif(card_addr_i = RCS) then
                        next_gen_state <= READOUT_CARD1;
                     elsif(card_addr_i = ALL_FBGA_CARDS) then
                        next_gen_state <= ADDR_CARD;
                     elsif(card_addr_i = ALL_CARDS) then
                        next_gen_state <= PS_CARD;
                     elsif(card_addr_i = PSC) then
                        next_gen_state <= PS_CARD;
                     elsif(card_addr_i = CC) then
                        next_gen_state <= CLOCK_CARD;
                     elsif(card_addr_i = AC) then
                        next_gen_state <= ADDR_CARD;
                     elsif(card_addr_i = RC1) then
                        next_gen_state <= READOUT_CARD1;
                     elsif(card_addr_i = RC2) then
                        next_gen_state <= READOUT_CARD2;
                     elsif(card_addr_i = RC3) then
                        next_gen_state <= READOUT_CARD3;
                     elsif(card_addr_i = RC4) then
                        next_gen_state <= READOUT_CARD4;
                     elsif(card_addr_i = BC1) then
                        next_gen_state <= BIAS_CARD1;
                     elsif(card_addr_i = BC2) then
                        next_gen_state <= BIAS_CARD2;
                     elsif(card_addr_i = BC3) then
                        next_gen_state <= BIAS_CARD3;
                     else
                        next_gen_state <= IDLE;  -- Catch all invalid card_id's with this statement
                     end if;
                  else
                     next_gen_state <= DONE;
                  end if;
               else
                  next_gen_state <= DONE;
               end if;
            else
               next_gen_state <= CLEANUP;
            end if;
         when DONE =>
            next_gen_state <= IDLE;
         when others =>
            next_gen_state <= IDLE;
      end case;
   end process;

   with card_addr_i(CARD_ADDR_WIDTH-1 downto 0) select
      cards_addressed <=
         0 when NO_CARDS,
         1 when PSC | CC | RC1 | RC2 | RC3 | RC4 | BC1 | BC2 | BC3 | AC,
         3 when BCS,
         4 when RCS,
         9 when ALL_FBGA_CARDS,
         10 when ALL_CARDS,
         0 when others; -- invalid card address

   -- The par_id checking is done in the cmd_translator block.
   -- Thus, here I can use the 'when others' case for something other than
   -- error checking, because the par_id that cmd_translator issues to cmd_queue
   -- is always valid.
   with par_id_i(7 downto 0) select
      uops_generated <=
         6 when RET_DAT_ADDR,
         5 when STATUS_ADDR,
         1 when others; -- all other m-ops generate one u-op

   num_uops <= uops_generated * cards_addressed;
   data_size_int <= conv_integer(data_size_i);
   size_uops <= num_uops * (2 + data_size_int);

   mop_rdy <= mop_rdy_i;

   gen_state_out: process(present_gen_state, par_id_i, card_addr_i) -- had new_card_addr_i
      begin
      case present_gen_state is
         when RESET =>
            insert_uop_rdy    <= '0';
            new_card_addr     <= card_addr_i(CQ_CARD_ADDR_BUS_WIDTH-1 downto 0);
            num_uops_inserted <= 0;
         when IDLE =>
            insert_uop_rdy    <= '0';
            new_card_addr     <= card_addr_i(CQ_CARD_ADDR_BUS_WIDTH-1 downto 0);
         when INSERT =>
            -- Add new u-ops to the queue
            insert_uop_rdy    <= '0';
            new_card_addr     <= card_addr_i(CQ_CARD_ADDR_BUS_WIDTH-1 downto 0);
            uop_counter       <= (others => '0');
            if(par_id_i(7 downto 0) = RET_DAT_ADDR) then
               new_par_id(7 downto 0) <= RET_DAT_ADDR;
            elsif(par_id_i(7 downto 0) = STATUS_ADDR) then
               new_par_id(7 downto 0) <= PSC_STATUS_ADDR;
            else
               new_par_id(7 downto 0) <= par_id_i(7 downto 0);
            end if;
         when PS_CARD | CLOCK_CARD | ADDR_CARD | READOUT_CARD1 | READOUT_CARD2 | READOUT_CARD3 | READOUT_CARD4 | BIAS_CARD1 | BIAS_CARD2 | BIAS_CARD3 =>
            insert_uop_rdy    <= '1';
            num_uops_inserted <= num_uops_inserted + 1;
            uop_counter       <= uop_counter + 1;
            if(present_gen_state = PS_CARD) then
               new_card_addr(CARD_ADDR_WIDTH-1 downto 0) <= PSC;
            elsif(present_gen_state = CLOCK_CARD) then
               new_card_addr(CARD_ADDR_WIDTH-1 downto 0) <= CC;
            elsif(present_gen_state = ADDR_CARD) then
               new_card_addr(CARD_ADDR_WIDTH-1 downto 0) <= AC;
            elsif(present_gen_state = READOUT_CARD1) then
               new_card_addr(CARD_ADDR_WIDTH-1 downto 0) <= RC1;
            elsif(present_gen_state = READOUT_CARD2) then
               new_card_addr(CARD_ADDR_WIDTH-1 downto 0) <= RC2;
            elsif(present_gen_state = READOUT_CARD3) then
               new_card_addr(CARD_ADDR_WIDTH-1 downto 0) <= RC3;
            elsif(present_gen_state = READOUT_CARD4) then
               new_card_addr(CARD_ADDR_WIDTH-1 downto 0) <= RC4;
            elsif(present_gen_state = BIAS_CARD1) then
               new_card_addr(CARD_ADDR_WIDTH-1 downto 0) <= BC1;
            elsif(present_gen_state = BIAS_CARD2) then
               new_card_addr(CARD_ADDR_WIDTH-1 downto 0) <= BC2;
            elsif(present_gen_state = BIAS_CARD3) then
               new_card_addr(CARD_ADDR_WIDTH-1 downto 0) <= BC3;
            end if;
         when CLEANUP =>
            insert_uop_rdy <= '0';
            new_card_addr  <= card_addr_i(CQ_CARD_ADDR_BUS_WIDTH-1 downto 0);
            if(par_id_i(7 downto 0) = RET_DAT_ADDR) then
               if(new_par_id(7 downto 0) = RET_DAT_ADDR) then
                  new_par_id(7 downto 0) <= PSC_STATUS_ADDR;
               elsif(new_par_id(7 downto 0) = PSC_STATUS_ADDR) then
                  new_par_id(7 downto 0) <= BIT_STATUS_ADDR;
               elsif(new_par_id(7 downto 0) = BIT_STATUS_ADDR) then
                  new_par_id(7 downto 0) <= FPGA_TEMP_ADDR;
               elsif(new_par_id(7 downto 0) = FPGA_TEMP_ADDR) then
                  new_par_id(7 downto 0) <= CARD_TEMP_ADDR;
               elsif(new_par_id(7 downto 0) = CARD_TEMP_ADDR) then
                  new_par_id(7 downto 0) <= CYC_OO_SYC_ADDR;
               elsif(new_par_id(7 downto 0) = CYC_OO_SYC_ADDR) then
                  new_par_id(7 downto 0) <= par_id_i(7 downto 0);
               end if;
            elsif(par_id_i(7 downto 0) = STATUS_ADDR) then
               if(new_par_id(7 downto 0) = PSC_STATUS_ADDR) then
                  new_par_id(7 downto 0) <= BIT_STATUS_ADDR;
               elsif(new_par_id(7 downto 0) = BIT_STATUS_ADDR) then
                  new_par_id(7 downto 0) <= FPGA_TEMP_ADDR;
               elsif(new_par_id(7 downto 0) = FPGA_TEMP_ADDR) then
                  new_par_id(7 downto 0) <= CARD_TEMP_ADDR;
               elsif(new_par_id(7 downto 0) = CARD_TEMP_ADDR) then
                  new_par_id(7 downto 0) <= CYC_OO_SYC_ADDR;
               elsif(new_par_id(7 downto 0) = CYC_OO_SYC_ADDR) then
                  new_par_id(7 downto 0) <= par_id_i(7 downto 0);
               end if;
            else
               new_par_id(7 downto 0) <= par_id_i(7 downto 0);
            end if;
         when DONE =>
            insert_uop_rdy    <= '0';
            new_card_addr     <= card_addr_i(CQ_CARD_ADDR_BUS_WIDTH-1 downto 0);
            num_uops_inserted <= 0;
         when others => -- Normal insertion
            insert_uop_rdy    <= '0';
            new_card_addr     <= card_addr_i(CQ_CARD_ADDR_BUS_WIDTH-1 downto 0);
      end case;
   end process;

   -- Send FSM:
   send_state_FF: process(clk_i, rst_i)
   begin
      if(rst_i = '1') then
         present_send_state <= RESET;
      elsif(clk_i'event and clk_i = '1') then
         present_send_state <= next_send_state;
      end if;
   end process send_state_FF;

   issue_sync       <= qa_sig(QUEUE_WIDTH-1 downto ISSUE_SYNC_END);
   timeout_sync     <= qa_sig(ISSUE_SYNC_END-1 downto TIMEOUT_SYNC_END);

   -- There should be enough time in the sync period following the timeout_sync of a m-op to get rid of all it's u-ops and still have time to issue the u-ops that need to be issued during that period
   -- That is why we don't check for a range here - just for the sync period that is the timeout
   -- This second conditions checks to see whether the instruction is in the black out period of the last valid sync pulse during which it can be issued.
   uop_send_expired <= '1' when (sync_count_slv = timeout_sync or
                                (sync_count_slv = timeout_sync - 1 and clk_count > START_OF_BLACKOUT)) else '0';

   send_state_NS: process(present_send_state, send_ptr, free_ptr, uop_send_expired, issue_sync, timeout_sync, sync_count_slv)
   begin
      case present_send_state is
         when RESET =>
            next_send_state <= LOAD;
         when LOAD =>
            -- If there is a u-op waiting to be issued, load it.  If not, idle
            if(send_ptr /= free_ptr) then
               if(uop_send_expired = '1') then
                  -- If the u-op has expired, it should be skipped
                  next_send_state <= NEXT_UOP;
               elsif(issue_sync < timeout_sync) then
                  -- Determine whether the current sync period is between the issue sync and the timeout sync.  If so, the u-op should be issued.
                  if(sync_count_slv >= issue_sync and sync_count_slv < timeout_sync) then
                     next_send_state <= HEADER_A;
                  else
                     next_send_state <= LOAD;
                  end if;
               -- The timeout_sync can have wrapped with respect to the issue_sync
               elsif(issue_sync > timeout_sync) then
                  if(sync_count_slv >= issue_sync or sync_count_slv < timeout_sync) then
                     next_send_state <= HEADER_A;
                  else
                     next_send_state <= LOAD;
                  end if;
               else
                  -- If the u-op is still good, but isn't supposed to be issued yet, stay in VERIFY
                  next_send_state <= LOAD;
               end if;
            elsif(send_ptr = free_ptr) then
               next_send_state <= LOAD;
            end if;
         when HEADER_A =>
            if(cmd_tx_done = '1' and crc_done = '1') then
               next_send_state <= HEADER_B;
            else
               next_send_state <= HEADER_A;
            end if;
         when HEADER_B =>
            if(cmd_tx_done = '1' and crc_done = '1') then
               if(there's data) then
                  next_send_state <= DATA;
               else
                  next_send_state <= CHECKSUM;
               end if;
            else
               next_send_state <= HEADER_B;
            end if;
         when DATA =>
            if(cmd_tx_done = '1' and crc_done = '1') then
               next_send_state <= CHECKSUM;
            else
               next_send_state <= DATA;
            end if;
         when CHECKSUM =>
            if(cmd_tx_done = '1') then
               next_send_state <= DONE;
            else
               next_send_state <= CHECKSUM;
            end if;
         when DONE =>
            next_send_state <= IDLE;
         when others =>
            next_send_state <= IDLE;
         when NEXT_UOP =>
            -- Skip to the next u-op
            next_send_state <= LOAD;
         when others =>
            next_send_state <= LOAD;
      end case;
   end process;

   rdaddress_a_sig <= send_ptr;

   send_state_out: process(present_send_state)
   begin
      case present_send_state is
         when RESET =>
            send_ptr   <= ADDR_ZERO;
         when LOAD =>
            tx_uop_rdy <= '0';
         when ISSUE =>
            -- All issue functionality may be contained in the Bus Backplane Packetization FSM
            tx_uop_rdy <= '1';
         when IDLE =>
            tx_uop_ack   <= '0';
            cmd_tx_start <= '0';
         when HEADER_A =>
            cmd_tx_start <= '1';
            -- Start of Command, 16 bits
            cmd_tx_dat(31 downto 16) <= x"AAAA";
            -- Size of Command, 16 bits
            cmd_tx_dat(15 downto  0) <= qa_sig(TIMEOUT_SYNC_END-1 downto DATA_SIZE_END);
         when HEADER_B =>
            cmd_tx_start <= '1';
            send_ptr   <= send_ptr + 1
--            cmd_tx_dat(31 downto 24) <= qa_sig(
--            cmd_tx_dat(23 downto 16) <=
--            cmd_tx_dat(15 downto  8) <=
--            cmd_tx_dat( 7 downto  0) <=
         when DATA =>
            cmd_tx_start <= '1';
            send_ptr   <= send_ptr + 1
         when CHECKSUM =>
            cmd_tx_start <= '1';
            send_ptr   <= send_ptr + 1
         when DONE =>
            cmd_tx_start <= '0';
         when others =>
            cmd_tx_start <= '0';
         when NEXT_UOP =>
            tx_uop_rdy <= '0';
            -- The send_ptr should be incremented in all situations, whether the u-op has expired or has been sent.
            send_ptr   <= send_ptr + 2 + qa_sig(DATA_SIZE_END+QUEUE_ADDR_WIDTH-1 downto DATA_SIZE_END);
         when others =>
            tx_uop_rdy <= '0';
      end case;
   end process;

   nfast_clk <= not clk_400mhz_i;
   n_clk <= not clk_i;
   sync_count_slv <= std_logic_vector(conv_unsigned(sync_count_int, 8));

end behav;

-- Bugs:
--x The insert FSM doesn't insert the first u-op in a sequence
--  I had to adjust the order that commands are issed over the bus backplane

--x The address card should be the last card that u-ops are issued to
--  There was a problem with what signals were on the sensitivity list.  For statements like i<=i+1, i should not appear in the sensitivity list

--x The generate FSM keeps on repeating the issue of u-ops to the AC
--  Solved by deasserting mop_rdy_o after mop_ack_i returned high

--x uops issued over the bus backplane should be issued in the following order: {for each uop(for each applicable card(issue uop))}
-- Done

--x the next_gen_state change occurs one clock cycle too late
--  added last_card_uop to the gen_NS fsm sensitivity list

--x last_card_uop count wrong.
-- removed last_card_uop becuase it is not used anymore.

--x new_card_addr should change one clock cycle earlier at the beginning of a sequence of u-ops issued
--  Done

--x the generate FSM cycles over two u-ops during a u-op transition
--  Done

--x uop_counter wraps at 31.  UOP_BUS_WIDTH is only bit bits wide.
--  UOP_BUS_WIDTH and MOP_BUS_WIDTH have been widened to 8 bits each.

--x I need to widen the RAM lines to 64 bits.
--  Done.

--x Change the handshaking protocol with the cmd_translator so that the ack signal is only asserted when the cmd_queue is done receiving a m-op.
--  This is already done by the Generate FSM

--x How do I convert and integer to a std_logic_vector
-- conv_std_logic_vector(name of vector, width of vector)
-- include ieee.std_logic_unsigned.all

--x Right now, determinig whether there is enough queue_space is calculated based on the number of u-ops that are inserted
-- it should actually be calculated based on the number of u-ops and how large each u-op is.

--x Change the clock frequency for the ram block and insertion FSM to clk_i instead of fast_clk_i
-- Done but not tested

--x Figure out how to take continuous data from the cmd_translator block
-- The insert FSM can take continuous data at the normal clock frequency
-- Once it is done, it asserts insert_uop_ack to let the generate FSM know that it's ready to receive the next u-op
-- While it is inserting the u-op and data, it asserts the inserting signal to all the queue-size FSM to alter the space available in the queue
-- To begin the continuous data stream, the insert FSM asserts the mop_ack_o line directly.

--x Slow down the insertion FSM so that everything works with the same clock.
-- To do this, I will have to implement a handshaking protocol to stall the generate FSM while the insert FSM is busy
-- The handshaking protocol between insert and generate FSMs has been implemented.
-- The handshaking signals used are insert_uop_rdy and insert_uop_ack
-- These signals are used exclusively for this purpose.

-- Send FSM must send out all relevant fields in the correct order, while creating a checksum on the fly

-- Check the sensitivity lists on the FSMs that I've been testing this morning.

-- Combine the packetization and send FSMs together, because they both need write access to send_ptr.

-- Write the supporting code in the send FSM for freeze_send.

-- Disable the CRC while the lvds_tx block finishes transmission.  
-- We are garunteed that the CRC block will finish calculating the checksum before the lvdsl_tx finishes tx'in the data

-- The 25Mhz LVDS clk should actually be 200 Mhz