-- Copyright (c) 2003 SCUBA-2 Project
--                  All Rights Reserved

--  THIS IS UNPUBLISHED PROPRIETARY SOURCE CODE OF THE SCUBA-2 Project
--  The copyright notice above does not evidence any
--  actual or intended publication of such source code.

--  SOURCE CODE IS PROVIDED "AS IS". ALL EXPRESS OR IMPLIED CONDITIONS,
--  REPRESENTATIONS, AND WARRANTIES, INCLUDING ANY IMPLIED WARRANT OF
--  MERCHANTABILITY, SATISFACTORY QUALITY, FITNESS FOR A PARTICULAR
--  PURPOSE, OR NON-INFRINGEMENT, ARE DISCLAIMED, EXCEPT TO THE EXTENT
--  THAT SUCH DISCLAIMERS ARE HELD TO BE LEGALLY INVALID.

-- For the purposes of this code the SCUBA-2 Project consists of the
-- following organisations.

-- UKATC, Royal Observatory, Blackford Hill Edinburgh EH9 3HJ
-- UBC,   University of British Columbia, Physics & Astronomy Department,
--        Vancouver BC, V6T 1Z1

-- frame_timing.vhd
--
-- <revision control keyword substitutions e.g. $Id: frame_timing.vhd,v 1.7 2004/05/17 22:33:06 mandana Exp $>
--
-- Project:		 SCUBA-2
-- Author:		 Bryce Burger
-- Organisation:	UBC
--
-- Description:
-- This implements the frame synchronization block for the AC, BC, RC.
--
-- Revision history:
-- <date $Date: 2004/05/17 22:33:06 $> - <text> - <initials $Author: mandana $>
-- $Log: frame_timing.vhd,v $
-- Revision 1.7  2004/05/17 22:33:06  mandana
-- changed counter output to integer
--
-- Revision 1.6  2004/04/16 23:30:21  mandana
-- fixed frame_rst
--
-- Revision 1.5  2004/04/16 21:58:05  bburger
-- bug fixes
--
-- Revision 1.4  2004/04/16 00:41:44  bburger
-- renamed some signals
--
-- Revision 1.3  2004/04/14 00:25:37  mandana
-- cleaned up extra signals
--
-- Revision 1.2  2004/04/03 01:05:37  bburger
-- Added a rst_on_next_sync_pulse register so that the master block doesn't have to assert that signal during the receipt of a sync, but anytime before
--
-- Revision 1.1  2004/04/02 01:13:13  bburger
-- New
--
--
------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

library sys_param;
use sys_param.frame_timing_pack.all;

library components;
use components.component_pack.all;

entity frame_timing is
   port(
      clk_i       : in std_logic;
      sync_i      : in std_logic;
      frame_rst_i : in std_logic;
      clk_count_o : out integer;
      clk_error_o : out std_logic_vector(31 downto 0)
   );
end frame_timing;

architecture beh of frame_timing is

   signal frame_rst : std_logic;
   signal clk_error : std_logic_vector(31 downto 0);
   signal counter_rst : std_logic;
   signal count : std_logic_vector(31 downto 0);
   signal count_int : integer;
   signal reg_rst : std_logic;
   type states is (WAIT_FRM_RST, WAIT_FOR_SYNC);
   
   signal current_state, next_state : states;
   
   begin
   cntr : counter
      generic map(MAX => END_OF_FRAME)
      port map(
         clk_i => clk_i,
         rst_i => counter_rst,
         ena_i => '1',
         load_i => '0',
         down_i => '0',
         count_i => 0,
         count_o => count_int
      );

   rstr : reg
      generic map(WIDTH => 32)
      port map(
         clk_i => sync_i,
         rst_i => reg_rst,
         ena_i => '1',
         reg_i  => count,
         reg_o => clk_error
      );

   count <= conv_std_logic_vector(count_int, 32);

   -- Inputs/Outputs
   clk_count_o <= count_int;
   clk_error_o <= clk_error;
   
-- CLOCKED FSMs
   state_FF: process(clk_i)
   begin
      if(clk_i'event and clk_i = '1') then
         current_state     <= next_state;
      end if;
   end process state_FF;

  state_NS: process(current_state, sync_i, frame_rst_i)
   begin
      case current_state is
         when WAIT_FRM_RST =>
            if frame_rst_i = '1' then
               next_state <= WAIT_FOR_SYNC;            
            end if;                  
         when WAIT_FOR_SYNC =>
            if (sync_i = '1') then
               next_state <= WAIT_FRM_RST;
            end if;
      end case;
   end process state_NS;
   
   counter_rst <= '1' when current_state = WAIT_FOR_SYNC and sync_i = '1' else '0';
   reg_rst     <= '1' when current_state = WAIT_FOR_SYNC and sync_i = '1' else '0';
   
end beh;