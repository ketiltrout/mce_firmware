-- megafunction wizard: %LPM_ADD_SUB%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: lpm_add_sub 

-- ============================================================
-- File Name: fsfb_calc_sub29.vhd
-- Megafunction Name(s):
-- 			lpm_add_sub
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 4.1 Build 208 09/10/2004 SP 2 SJ Full Version
-- ************************************************************


--Copyright (C) 1991-2004 Altera Corporation
--Any  megafunction  design,  and related netlist (encrypted  or  decrypted),
--support information,  device programming or simulation file,  and any other
--associated  documentation or information  provided by  Altera  or a partner
--under  Altera's   Megafunction   Partnership   Program  may  be  used  only
--to program  PLD  devices (but not masked  PLD  devices) from  Altera.   Any
--other  use  of such  megafunction  design,  netlist,  support  information,
--device programming or simulation file,  or any other  related documentation
--or information  is prohibited  for  any  other purpose,  including, but not
--limited to  modification,  reverse engineering,  de-compiling, or use  with
--any other  silicon devices,  unless such use is  explicitly  licensed under
--a separate agreement with  Altera  or a megafunction partner.  Title to the
--intellectual property,  including patents,  copyrights,  trademarks,  trade
--secrets,  or maskworks,  embodied in any such megafunction design, netlist,
--support  information,  device programming or simulation file,  or any other
--related documentation or information provided by  Altera  or a megafunction
--partner, remains with Altera, the megafunction partner, or their respective
--licensors. No other licenses, including any licenses needed under any third
--party's intellectual property, are provided herein.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY fsfb_calc_sub29 IS
	PORT
	(
		dataa		: IN STD_LOGIC_VECTOR (28 DOWNTO 0);
		datab		: IN STD_LOGIC_VECTOR (28 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (28 DOWNTO 0)
	);
END fsfb_calc_sub29;


ARCHITECTURE SYN OF fsfb_calc_sub29 IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (28 DOWNTO 0);



	COMPONENT lpm_add_sub
	GENERIC (
		lpm_width		: NATURAL;
		lpm_direction		: STRING;
		lpm_type		: STRING;
		lpm_hint		: STRING
	);
	PORT (
			dataa	: IN STD_LOGIC_VECTOR (28 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (28 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (28 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(28 DOWNTO 0);

	lpm_add_sub_component : lpm_add_sub
	GENERIC MAP (
		lpm_width => 29,
		lpm_direction => "SUB",
		lpm_type => "LPM_ADD_SUB",
		lpm_hint => "ONE_INPUT_IS_CONSTANT=NO,CIN_USED=NO"
	)
	PORT MAP (
		dataa => dataa,
		datab => datab,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: nBit NUMERIC "29"
-- Retrieval info: PRIVATE: Function NUMERIC "1"
-- Retrieval info: PRIVATE: RadixA NUMERIC "10"
-- Retrieval info: PRIVATE: RadixB NUMERIC "10"
-- Retrieval info: PRIVATE: WhichConstant NUMERIC "0"
-- Retrieval info: PRIVATE: ConstantA NUMERIC "0"
-- Retrieval info: PRIVATE: ConstantB NUMERIC "0"
-- Retrieval info: PRIVATE: ValidCtA NUMERIC "0"
-- Retrieval info: PRIVATE: ValidCtB NUMERIC "0"
-- Retrieval info: PRIVATE: CarryIn NUMERIC "0"
-- Retrieval info: PRIVATE: CarryOut NUMERIC "0"
-- Retrieval info: PRIVATE: Overflow NUMERIC "0"
-- Retrieval info: PRIVATE: Latency NUMERIC "0"
-- Retrieval info: PRIVATE: aclr NUMERIC "0"
-- Retrieval info: PRIVATE: clken NUMERIC "0"
-- Retrieval info: PRIVATE: LPM_PIPELINE NUMERIC "0"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "29"
-- Retrieval info: CONSTANT: LPM_DIRECTION STRING "SUB"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_ADD_SUB"
-- Retrieval info: CONSTANT: LPM_HINT STRING "ONE_INPUT_IS_CONSTANT=NO,CIN_USED=NO"
-- Retrieval info: USED_PORT: result 0 0 29 0 OUTPUT NODEFVAL result[28..0]
-- Retrieval info: USED_PORT: dataa 0 0 29 0 INPUT NODEFVAL dataa[28..0]
-- Retrieval info: USED_PORT: datab 0 0 29 0 INPUT NODEFVAL datab[28..0]
-- Retrieval info: CONNECT: result 0 0 29 0 @result 0 0 29 0
-- Retrieval info: CONNECT: @dataa 0 0 29 0 dataa 0 0 29 0
-- Retrieval info: CONNECT: @datab 0 0 29 0 datab 0 0 29 0
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL fsfb_calc_sub29.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fsfb_calc_sub29.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fsfb_calc_sub29.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fsfb_calc_sub29.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fsfb_calc_sub29_inst.vhd FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fsfb_calc_sub29_waveforms.html FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fsfb_calc_sub29_wave*.jpg FALSE
