-- Copyright (c) 2003 SCUBA-2 Project
--                  All Rights Reserved
--
--  THIS IS UNPUBLISHED PROPRIETARY SOURCE CODE OF THE SCUBA-2 Project
--  The copyright notice above does not evidence any
--  actual or intended publication of such source code.
--
--  SOURCE CODE IS PROVIDED "AS IS". ALL EXPRESS OR IMPLIED CONDITIONS,
--  REPRESENTATIONS, AND WARRANTIES, INCLUDING ANY IMPLIED WARRANT OF
--  MERCHANTABILITY, SATISFACTORY QUALITY, FITNESS FOR A PARTICULAR
--  PURPOSE, OR NON-INFRINGEMENT, ARE DISCLAIMED, EXCEPT TO THE EXTENT
--  THAT SUCH DISCLAIMERS ARE HELD TO BE LEGALLY INVALID.
--
-- For the purposes of this code the SCUBA-2 Project consists of the
-- following organisations.
--
-- UKATC, Royal Observatory, Blackford Hill Edinburgh EH9 3HJ
-- UBC,   University of British Columbia, Physics & Astronomy Department,
--        Vancouver BC, V6T 1Z1
--
--
-- p_banks_admin.vhd
--
-- Project:	  SCUBA-2
-- Author:        Mohsen Nahvi
-- Organisation:  UBC
--
-- Description:
-- 
-- This block instantiates the P memory RAMs for each 8 channel of the
-- flux_loop_ctrl.  The memory banks are registered both at the inputs and the
-- outputs.  Therefore, a write cycle is complete on the next rising edge
-- of the clock after the address is valid.  However, a read cycle is only
-- complete after two clock cycles after the address is valid. (NOTE: that the
-- data can be read on the third clock rising edge)
--
-- Two control signals are also generated.
-- 1. The first one is the write enable signal for each memory bank.  These
-- signals are simply the we_i when the addr_i is equal to the address of that
-- memory bank.
-- 2. The second control signal is the ack_o.  This signal is generated
-- separtely for each of the write or read cycle.  A behavioural code is used
-- for simplicity where the idea is to generate the ack_o every other clock
-- cycles during a write and every two other clock cycles during a read.
--
-- Ports:
-- #clk_50_i: Golbal signal
-- #rst_i: Global signal
-- #p_dat_ch0_o: P Data for flux_loop_ctrl channel0
-- #p_addr_ch0_i: Read address from flux_loop_ctrl channle0
-- #### Similarly for ch1 to ch7
-- #dat_i: Data in from Dispatch
-- #addr_i: Address from Dispatch showing the address of memory banks. This is
-- kept constant during a read or write cycle.
-- #tga_i: Address Tag from Dispatch.  This is incremented during a read or
-- write cycle.  Therefore, it is used as an index to the location in the
-- memory bank
-- #we_i: Write Enable input from Dispatch
-- #stb_i: Strobe signal from Dispatch.  Indicates if an address is valid or
-- not. See Wishbone manul page 54 and 57.  
-- #cyc_i: Input from Dispatch indicating a read or write cycle is in progress
-- #qa_p_bank_o: A MUX output of all the qa output of the memory banks for P 
-- #ack_p_bank_o: A logical OR function of acknowledge signals for read or
-- write cycles of each memory bank
--
--
--
-- Revision history:
-- 
-- $Log: p_banks_admin.vhd,v $
-- Revision 1.1  2004/11/20 01:22:02  mohsen
-- Initial release
--
--
--
------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

library sys_param;
use sys_param.command_pack.all;
use sys_param.wishbone_pack.all;

library work;

-- Call Parent Library
use work.wbs_fb_data_pack.all;
use work.flux_loop_pack.all;



entity p_banks_admin is
  
  port (

    -- Global signals
    clk_50_i                : in std_logic;
    rst_i                   : in std_logic;


    -- Flux_Loop_Ctrl Channel Interface
    p_dat_ch0_o             : out std_logic_vector(WB_DATA_WIDTH-1 downto 0);   
    p_addr_ch0_i            : in  std_logic_vector(PIDZ_ADDR_WIDTH-1 downto 0);   
    p_dat_ch1_o             : out std_logic_vector(WB_DATA_WIDTH-1 downto 0);   
    p_addr_ch1_i            : in  std_logic_vector(PIDZ_ADDR_WIDTH-1 downto 0);   
    p_dat_ch2_o             : out std_logic_vector(WB_DATA_WIDTH-1 downto 0);   
    p_addr_ch2_i            : in  std_logic_vector(PIDZ_ADDR_WIDTH-1 downto 0);   
    p_dat_ch3_o             : out std_logic_vector(WB_DATA_WIDTH-1 downto 0);   
    p_addr_ch3_i            : in  std_logic_vector(PIDZ_ADDR_WIDTH-1 downto 0);   
    p_dat_ch4_o             : out std_logic_vector(WB_DATA_WIDTH-1 downto 0);   
    p_addr_ch4_i            : in  std_logic_vector(PIDZ_ADDR_WIDTH-1 downto 0);   
    p_dat_ch5_o             : out std_logic_vector(WB_DATA_WIDTH-1 downto 0);   
    p_addr_ch5_i            : in  std_logic_vector(PIDZ_ADDR_WIDTH-1 downto 0);   
    p_dat_ch6_o             : out std_logic_vector(WB_DATA_WIDTH-1 downto 0);   
    p_addr_ch6_i            : in  std_logic_vector(PIDZ_ADDR_WIDTH-1 downto 0);   
    p_dat_ch7_o             : out std_logic_vector(WB_DATA_WIDTH-1 downto 0);   
    p_addr_ch7_i            : in  std_logic_vector(PIDZ_ADDR_WIDTH-1 downto 0);
    

    -- signals to/from dispatch  (wishbone interface)
    dat_i                   : in  std_logic_vector(WB_DATA_WIDTH-1 downto 0);       -- wishbone data in
    addr_i                  : in  std_logic_vector(WB_ADDR_WIDTH-1 downto 0);       -- wishbone address in
    tga_i                   : in  std_logic_vector(WB_TAG_ADDR_WIDTH-1 downto 0);   -- Address Tag
    we_i                    : in  std_logic;                                        -- write//read enable
    stb_i                   : in  std_logic;                                        -- strobe 
    cyc_i                   : in  std_logic;                                        -- cycle
    --dat_o                   : out std_logic_vector(WB_DATA_WIDTH-1 downto 0);       -- data out
    --ack_o                   : out std_logic;                                        -- acknowledge out
    
    
    -- Interface intended for dispatch
    qa_p_bank_o             : out std_logic_vector(WB_DATA_WIDTH-1 downto 0);
    ack_p_bank_o            : out std_logic);
  

end p_banks_admin;



architecture rtl of p_banks_admin is

  -----------------------------------------------------------------------------
  -- Signals from P Banks
  -----------------------------------------------------------------------------
  signal qa_p_bank_ch0 : std_logic_vector(WB_DATA_WIDTH-1 downto 0);
  signal qa_p_bank_ch1 : std_logic_vector(WB_DATA_WIDTH-1 downto 0);
  signal qa_p_bank_ch2 : std_logic_vector(WB_DATA_WIDTH-1 downto 0);
  signal qa_p_bank_ch3 : std_logic_vector(WB_DATA_WIDTH-1 downto 0);
  signal qa_p_bank_ch4 : std_logic_vector(WB_DATA_WIDTH-1 downto 0);
  signal qa_p_bank_ch5 : std_logic_vector(WB_DATA_WIDTH-1 downto 0);
  signal qa_p_bank_ch6 : std_logic_vector(WB_DATA_WIDTH-1 downto 0);
  signal qa_p_bank_ch7 : std_logic_vector(WB_DATA_WIDTH-1 downto 0);

  
  -----------------------------------------------------------------------------
  -- Signals from P Controller
  -----------------------------------------------------------------------------
  signal wren_p_bank_ch0  : std_logic;
  signal wren_p_bank_ch1  : std_logic;
  signal wren_p_bank_ch2  : std_logic;
  signal wren_p_bank_ch3  : std_logic;
  signal wren_p_bank_ch4  : std_logic;
  signal wren_p_bank_ch5  : std_logic;
  signal wren_p_bank_ch6  : std_logic;
  signal wren_p_bank_ch7  : std_logic;
  signal ack_read_p_bank  : std_logic;
  signal ack_write_p_bank : std_logic;


  
begin  -- rtl


  -----------------------------------------------------------------------------
  -- Instantiation of P Banks
  -----------------------------------------------------------------------------

  i_p_bank_ch0 : wbs_fb_storage
    port map (
    data        => dat_i,                             -- from dispatch
    wraddress   => tga_i(PIDZ_ADDR_WIDTH-1 downto 0), -- from dispatch
    rdaddress_a => tga_i(PIDZ_ADDR_WIDTH-1 downto 0), -- from dispatch
    rdaddress_b => p_addr_ch0_i,                      -- from flux_loop_ctrl ch0
    wren        => wren_p_bank_ch0,                   -- from controller
    clock       => clk_50_i,                          -- global input
    qa          => qa_p_bank_ch0,                     -- to output intended for dispatch
    qb          => p_dat_ch0_o);                      -- to flux_loop_ctrl ch0
  

  i_p_bank_ch1 : wbs_fb_storage
    port map (
    data        => dat_i,                             -- from dispatch
    wraddress   => tga_i(PIDZ_ADDR_WIDTH-1 downto 0), -- from dispatch
    rdaddress_a => tga_i(PIDZ_ADDR_WIDTH-1 downto 0), -- from dispatch
    rdaddress_b => p_addr_ch1_i,                      -- from flux_loop_ctrl ch1
    wren        => wren_p_bank_ch1,                   -- from controller
    clock       => clk_50_i,                          -- global input
    qa          => qa_p_bank_ch1,                     -- to output intended for dispatch
    qb          => p_dat_ch1_o);                      -- to flux_loop_ctrl ch1

  
  i_p_bank_ch2 : wbs_fb_storage
    port map (
    data        => dat_i,                             -- from dispatch
    wraddress   => tga_i(PIDZ_ADDR_WIDTH-1 downto 0), -- from dispatch
    rdaddress_a => tga_i(PIDZ_ADDR_WIDTH-1 downto 0), -- from dispatch
    rdaddress_b => p_addr_ch2_i,                      -- from flux_loop_ctrl ch2
    wren        => wren_p_bank_ch2,                   -- from controller
    clock       => clk_50_i,                          -- global input
    qa          => qa_p_bank_ch2,                     -- to output intended for dispatch
    qb          => p_dat_ch2_o);                      -- to flux_loop_ctrl ch2


  i_p_bank_ch3 : wbs_fb_storage
    port map (
    data        => dat_i,                             -- from dispatch
    wraddress   => tga_i(PIDZ_ADDR_WIDTH-1 downto 0), -- from dispatch
    rdaddress_a => tga_i(PIDZ_ADDR_WIDTH-1 downto 0), -- from dispatch
    rdaddress_b => p_addr_ch3_i,                      -- from flux_loop_ctrl ch3
    wren        => wren_p_bank_ch3,                   -- from controller
    clock       => clk_50_i,                          -- global input
    qa          => qa_p_bank_ch3,                     -- to output intended for dispatch
    qb          => p_dat_ch3_o);                      -- to flux_loop_ctrl ch3


  i_p_bank_ch4 : wbs_fb_storage
    port map (
    data        => dat_i,                             -- from dispatch
    wraddress   => tga_i(PIDZ_ADDR_WIDTH-1 downto 0), -- from dispatch
    rdaddress_a => tga_i(PIDZ_ADDR_WIDTH-1 downto 0), -- from dispatch
    rdaddress_b => p_addr_ch4_i,                      -- from flux_loop_ctrl ch4
    wren        => wren_p_bank_ch4,                   -- from controller
    clock       => clk_50_i,                          -- global input
    qa          => qa_p_bank_ch4,                     -- to output intended for dispatch
    qb          => p_dat_ch4_o);                      -- to flux_loop_ctrl ch4


  i_p_bank_ch5 : wbs_fb_storage
    port map (
    data        => dat_i,                             -- from dispatch
    wraddress   => tga_i(PIDZ_ADDR_WIDTH-1 downto 0), -- from dispatch
    rdaddress_a => tga_i(PIDZ_ADDR_WIDTH-1 downto 0), -- from dispatch
    rdaddress_b => p_addr_ch5_i,                      -- from flux_loop_ctrl ch5
    wren        => wren_p_bank_ch5,                   -- from controller
    clock       => clk_50_i,                          -- global input
    qa          => qa_p_bank_ch5,                     -- to output intended for dispatch
    qb          => p_dat_ch5_o);                      -- to flux_loop_ctrl ch5
  

  i_p_bank_ch6 : wbs_fb_storage
    port map (
    data        => dat_i,                             -- from dispatch
    wraddress   => tga_i(PIDZ_ADDR_WIDTH-1 downto 0), -- from dispatch
    rdaddress_a => tga_i(PIDZ_ADDR_WIDTH-1 downto 0), -- from dispatch
    rdaddress_b => p_addr_ch6_i,                      -- from flux_loop_ctrl ch6
    wren        => wren_p_bank_ch6,                   -- from controller
    clock       => clk_50_i,                          -- global input
    qa          => qa_p_bank_ch6,                     -- to output intended for dispatch
    qb          => p_dat_ch6_o);                      -- to flux_loop_ctrl ch6


  i_p_bank_ch7 : wbs_fb_storage
    port map (
    data        => dat_i,                             -- from dispatch
    wraddress   => tga_i(PIDZ_ADDR_WIDTH-1 downto 0), -- from dispatch
    rdaddress_a => tga_i(PIDZ_ADDR_WIDTH-1 downto 0), -- from dispatch
    rdaddress_b => p_addr_ch7_i,                      -- from flux_loop_ctrl ch7
    wren        => wren_p_bank_ch7,                   -- from controller
    clock       => clk_50_i,                          -- global input
    qa          => qa_p_bank_ch7,                     -- to output intended for dispatch
    qb          => p_dat_ch7_o);                      -- to flux_loop_ctrl ch7


  
  -----------------------------------------------------------------------------
  -- Controller for P Banks:
  -- 
  -- 1. Write Enable signals for each bank is equal to the dispatch we_i when
  -- the address from dispatch, addr_i, is equla to that bank's address
  --
  -- 2. Acknowledge signals are different for Write or Read cycle.
  -- 
  -- 2.1 Write Cycle:
  -- The acknowlege signal is asserted for one clock cycle on the first clock
  -- rising edge after seeing the stb_i, and repeats every other clock as long
  -- as stb_i is high.  Note that stb_i remains high if slave is asserting wait
  -- states, like our case here.  However, if the master is inserting a wait
  -- state, stb_i goes low on seeing acknowlege signal and comes back high when
  -- the master is ready.  We implement the Write acknowlege using a
  -- behavioural code.
  --
  -- 2.2 Read Cycle:
  -- The acknowlege signal is asserted for one clock cycle on the second clcok
  -- rising edge after seeing the stb_i, and repeats every 2 clock cycles as
  -- long as stb_i is high.  This is necessary as we use memory with registered
  -- outputs, and, thus, there are two clock cycles delay for the output to be
  -- ready on each read value.  We implement the Read acknowlege using a
  -- behavioural code.
  -----------------------------------------------------------------------------

  -----------------------------------------------------------------------------
  -- Write Enable Signals
  wren_p_bank_ch0 <=
    we_i when addr_i=GAINP0_ADDR else
    '0';
  
  wren_p_bank_ch1 <=
    we_i when addr_i=GAINP1_ADDR else
    '0';

  wren_p_bank_ch2 <=
    we_i when addr_i=GAINP2_ADDR else
    '0';

  wren_p_bank_ch3 <=
    we_i when addr_i=GAINP3_ADDR else
    '0';

  wren_p_bank_ch4 <=
    we_i when addr_i=GAINP4_ADDR else
    '0';

  wren_p_bank_ch5 <=
    we_i when addr_i=GAINP5_ADDR else
    '0';

  wren_p_bank_ch6 <=
    we_i when addr_i=GAINP6_ADDR else
    '0';

  wren_p_bank_ch7 <=
    we_i when addr_i=GAINP7_ADDR else
    '0';

  -----------------------------------------------------------------------------
  -- Acknowlege signals
  i_gen_ack: process (clk_50_i, rst_i)
    
    variable count : integer;           -- counts number of clock cycles passed
    
  begin  -- process i_gen_ack
    if rst_i = '1' then                 -- asynchronous reset (active high)
      ack_read_p_bank  <= '0';
      ack_write_p_bank <= '0';
      count:=0;
      
      
    elsif clk_50_i'event and clk_50_i = '1' then  -- rising clock edge
      
      -- Write Acknowledge
      if (we_i='1') and ((addr_i= GAINP0_ADDR) or
                         (addr_i= GAINP1_ADDR) or
                         (addr_i= GAINP2_ADDR) or
                         (addr_i= GAINP3_ADDR) or
                         (addr_i= GAINP4_ADDR) or
                         (addr_i= GAINP5_ADDR) or
                         (addr_i= GAINP6_ADDR) or
                         (addr_i= GAINP7_ADDR)) then
        
        if (stb_i='1') and (ack_write_p_bank='0') then
          ack_write_p_bank <= '1';
        else
          ack_write_p_bank <= '0';
        end if;
      else
        ack_write_p_bank <= '0';
      end if;

      
      -- Read Acknowledge
      if (we_i='0') and ((addr_i= GAINP0_ADDR) or
                         (addr_i= GAINP1_ADDR) or
                         (addr_i= GAINP2_ADDR) or
                         (addr_i= GAINP3_ADDR) or
                         (addr_i= GAINP4_ADDR) or
                         (addr_i= GAINP5_ADDR) or
                         (addr_i= GAINP6_ADDR) or
                         (addr_i= GAINP7_ADDR)) then
        
        if (stb_i='1') and (ack_read_p_bank='0') then
          count:=count+1;
          if count=2 then
            ack_read_p_bank <= '1';
            count:=0;
          end if;
        else
          ack_read_p_bank <= '0';
        end if;
        
        
      else
        ack_read_p_bank <= '0';
        
      end if;

      
    end if;
  end process i_gen_ack;



  
  -----------------------------------------------------------------------------
  -- Output MUX to Dispatch:
  -- 
  -- 1. addr_i selects which bank is sending its output to the dispatch.  The
  -- defulat connection is to ch0.
  --
  -- 2. Acknowlege is ORing of the write and read cycle
  -----------------------------------------------------------------------------

  ack_p_bank_o <= ack_write_p_bank or ack_read_p_bank;

  with addr_i select
    qa_p_bank_o <=
    qa_p_bank_ch0 when GAINP0_ADDR,
    qa_p_bank_ch1 when GAINP1_ADDR,
    qa_p_bank_ch2 when GAINP2_ADDR,
    qa_p_bank_ch3 when GAINP3_ADDR,
    qa_p_bank_ch4 when GAINP4_ADDR,
    qa_p_bank_ch5 when GAINP5_ADDR,
    qa_p_bank_ch6 when GAINP6_ADDR,
    qa_p_bank_ch7 when GAINP7_ADDR,
    qa_p_bank_ch0 when others;        -- default to ch0

  
  
end rtl;
