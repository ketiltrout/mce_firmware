-- Copyright (c) 2003 SCUBA-2 Project
--                  All Rights Reserved

--  THIS IS UNPUBLISHED PROPRIETARY SOURCE CODE OF THE SCUBA-2 Project
--  The copyright notice above does not evidence any
--  actual or intended publication of such source code.

--  SOURCE CODE IS PROVIDED "AS IS". ALL EXPRESS OR IMPLIED CONDITIONS,
--  REPRESENTATIONS, AND WARRANTIES, INCLUDING ANY IMPLIED WARRANT OF
--  MERCHANTABILITY, SATISFACTORY QUALITY, FITNESS FOR A PARTICULAR
--  PURPOSE, OR NON-INFRINGEMENT, ARE DISCLAIMED, EXCEPT TO THE EXTENT
--  THAT SUCH DISCLAIMERS ARE HELD TO BE LEGALLY INVALID.

-- For the purposes of this code the SCUBA-2 Project consists of the
-- following organisations.

-- UKATC, Royal Observatory, Blackford Hill Edinburgh EH9 3HJ
-- UBC,   University of British Columbia, Physics & Astronomy Department,
--        Vancouver BC, V6T 1Z1

-- 
--
-- <revision control keyword substitutions e.g. $Id: fibre_rx_fifo.vhd,v 1.4 2004/11/24 01:15:52 bench2 Exp $>
--
-- Project:       SCUBA-2
-- Author:        David Atkinson
--               
-- Organisation:  UK ATC
--
-- Description: Fibre optic Receive FIFO.   Bytes of data from the hotlink 
-- receiver are written to this FIFO.  Writing to this block
-- is controlled by rx_control block (with signals from HOTLINK receiver).
-- 
-- The FIFO needs to be deep enought to buffer one MCE command (at least 256 bytes)
--
-- Revision history:
-- 1st March 2004   - Initial version      - DA
-- 
-- <date $Date: 2004/11/24 01:15:52 $> -     <text>      - <initials $Author: bench2 $>
--
-- $Log: fibre_rx_fifo.vhd,v $
-- Revision 1.4  2004/11/24 01:15:52  bench2
-- Greg: Broke apart issue reply and created pack files for all of its sub-components
--
-- Revision 1.3  2004/10/11 13:31:27  dca
-- Now instantiates synchronous FIFO megafunction
--
-----------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
--use ieee.numeric_std.all;

library work;
use work.issue_reply_pack.all;
use work.fibre_rx_pack.all;

library components;
use components.component_pack.all;

--library sys_param;
--use sys_param.command_pack.all;

entity fibre_rx_fifo is
--   generic(addr_size : Positive);                                          -- use this if instantiating async fifo
   port( 
      clk_i        : in     std_logic;                                          -- global clock
      rst_i        : in     std_logic;                                          -- global reset
           
      fibre_clkr_i : in     std_logic;                                          -- CKR from hotlink receiver 
      rx_fr_i      : in     std_logic;                                          -- fifo read request
      rx_fw_i      : in     std_logic;                                          -- fifo write request
      rx_data_i    : in     std_logic_vector (RX_FIFO_DATA_WIDTH-1 downto 0);   -- fifo data input
      rx_fe_o      : out    std_logic;                                          -- fifo empty flag
      rx_ff_o      : out    std_logic;                                          -- fifo full flagg
      rxd_o        : out    std_logic_vector (RX_FIFO_DATA_WIDTH-1 downto 0)    -- fifo data output
   );

end fibre_rx_fifo ;


architecture rtl of fibre_rx_fifo is
   component sync_fifo_rx
	PORT
	(
		data		: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		wrreq		: IN STD_LOGIC ;
		rdreq		: IN STD_LOGIC ;
		rdclk		: IN STD_LOGIC ;
		wrclk		: IN STD_LOGIC ;
		aclr		: IN STD_LOGIC  := '0';
		q		: OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		rdempty		: OUT STD_LOGIC ;
		wrfull		: OUT STD_LOGIC 
	);
   END component;

begin
 
   -- instantiate asynchronous FIFO
   -- Instance port mappings.
--   AFIFO : async_fifo
--      generic map(addr_size => addr_size)
--     port map(
--         rst_i    => rst_i,
--         read_i   => rx_fr_i,
--         write_i  => rx_fw_i,
--         d_i      => rx_data_i,
--         empty_o  => rx_fe_o,
--         full_o   => rx_ff_o,
--        q_o      => rxd_o
--      );
  
  
   -- instantiate synchronous fifo
    
   SFIFO : sync_fifo_rx
   port map(
      data     => rx_data_i,
      wrreq    => rx_fw_i,
      rdreq    => rx_fr_i,
      rdclk    => clk_i, 
      wrclk    => fibre_clkr_i,
      aclr     => rst_i,    
      q     => rxd_o, 
      rdempty     => rx_fe_o, 
      wrfull      => rx_ff_o
      );  
  
end rtl;
